module riscv_decode (
    input logic [31:0] data,
    output logic ADD,
    output logic ADDI,
    output logic AND,
    output logic ANDI,
    output logic AUIPC,
    output logic BEQ,
    output logic BGE,
    output logic BGEU,
    output logic BLT,
    output logic BLTU,
    output logic BNE,
    output logic C_ADD,
    output logic C_ADDI,
    output logic C_ADDI16SP,
    output logic C_ADDI4SPN,
    output logic C_AND,
    output logic C_ANDI,
    output logic C_BEQZ,
    output logic C_BNEZ,
    output logic C_EBREAK,
    output logic C_J,
    output logic C_JAL,
    output logic C_JALR,
    output logic C_JR,
    output logic C_LI,
    output logic C_LUI,
    output logic C_LW,
    output logic C_LWSP,
    output logic C_MV,
    output logic C_NOP,
    output logic C_OR,
    output logic C_SUB,
    output logic C_SW,
    output logic C_SWSP,
    output logic C_XOR,
    output logic DIV,
    output logic DIVU,
    output logic EBREAK,
    output logic ECALL,
    output logic FENCE,
    output logic JAL,
    output logic JALR,
    output logic LB,
    output logic LBU,
    output logic LH,
    output logic LHU,
    output logic LUI,
    output logic LW,
    output logic MUL,
    output logic MULH,
    output logic MULHSU,
    output logic MULHU,
    output logic OR,
    output logic ORI,
    output logic REM,
    output logic REMU,
    output logic SB,
    output logic SH,
    output logic SLL,
    output logic SLT,
    output logic SLTI,
    output logic SLTIU,
    output logic SLTU,
    output logic SRA,
    output logic SRL,
    output logic SUB,
    output logic SW,
    output logic XOR,
    output logic XORI,
    output logic defined,
    output logic compressed,
    output logic bimm12hi,
    output logic bimm12lo,
    output logic c_bimm9hi,
    output logic c_bimm9lo,
    output logic c_imm12,
    output logic c_imm6hi,
    output logic c_imm6lo,
    output logic c_nzimm10hi,
    output logic c_nzimm10lo,
    output logic c_nzimm18hi,
    output logic c_nzimm18lo,
    output logic c_nzimm6hi,
    output logic c_nzimm6lo,
    output logic c_nzuimm10,
    output logic c_rs2,
    output logic c_uimm7hi,
    output logic c_uimm7lo,
    output logic c_uimm8sp_s,
    output logic c_uimm8sphi,
    output logic c_uimm8splo,
    output logic fm,
    output logic imm12,
    output logic imm12hi,
    output logic imm12lo,
    output logic imm20,
    output logic jimm20,
    output logic pred,
    output logic rd,
    output logic rd_p,
    output logic rd_rs1,
    output logic rd_rs1_p,
    output logic rs1,
    output logic rs1_p,
    output logic rs2,
    output logic rs2_p,
    output logic succ
);
   //ADD
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????000?????0110011: ADD = '1;
         default: ADD = '0;
      endcase
   end
   //ADDI
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????0010011: ADDI = '1;
         default: ADDI = '0;
      endcase
   end
   //AND
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????111?????0110011: AND = '1;
         default: AND = '0;
      endcase
   end
   //ANDI
   always_comb begin
      casez (data[31:0])
         32'b?????????????????111?????0010011: ANDI = '1;
         default: ANDI = '0;
      endcase
   end
   //AUIPC
   always_comb begin
      casez (data[31:0])
         32'b?????????????????????????0010111: AUIPC = '1;
         default: AUIPC = '0;
      endcase
   end
   //BEQ
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????1100011: BEQ = '1;
         default: BEQ = '0;
      endcase
   end
   //BGE
   always_comb begin
      casez (data[31:0])
         32'b?????????????????101?????1100011: BGE = '1;
         default: BGE = '0;
      endcase
   end
   //BGEU
   always_comb begin
      casez (data[31:0])
         32'b?????????????????111?????1100011: BGEU = '1;
         default: BGEU = '0;
      endcase
   end
   //BLT
   always_comb begin
      casez (data[31:0])
         32'b?????????????????100?????1100011: BLT = '1;
         default: BLT = '0;
      endcase
   end
   //BLTU
   always_comb begin
      casez (data[31:0])
         32'b?????????????????110?????1100011: BLTU = '1;
         default: BLTU = '0;
      endcase
   end
   //BNE
   always_comb begin
      casez (data[31:0])
         32'b?????????????????001?????1100011: BNE = '1;
         default: BNE = '0;
      endcase
   end
   //C_ADD
   always_comb begin
      casez (data[31:0])
         32'b????????????????1001????????1?10: C_ADD = '1;
         32'b????????????????1001??????1???10: C_ADD = '1;
         32'b????????????????1001???????1??10: C_ADD = '1;
         32'b????????????????1001?????1????10: C_ADD = '1;
         32'b????????????????1001?????????110: C_ADD = '1;
         default: C_ADD = '0;
      endcase
   end
   //C_ADDI
   always_comb begin
      casez (data[31:0])
         32'b????????????????000?1?????????01: C_ADDI = '1;
         32'b????????????????000??1????????01: C_ADDI = '1;
         32'b????????????????000?????1?????01: C_ADDI = '1;
         32'b????????????????000???1???????01: C_ADDI = '1;
         32'b????????????????000????1??????01: C_ADDI = '1;
         default: C_ADDI = '0;
      endcase
   end
   //C_ADDI16SP
   always_comb begin
      casez (data[31:0])
         32'b????????????????011?00010?????01: C_ADDI16SP = '1;
         default: C_ADDI16SP = '0;
      endcase
   end
   //C_ADDI4SPN
   always_comb begin
      casez (data[31:0])
         32'b????????????????000???????????00: C_ADDI4SPN = '1;
         default: C_ADDI4SPN = '0;
      endcase
   end
   //C_AND
   always_comb begin
      casez (data[31:0])
         32'b????????????????100011???11???01: C_AND = '1;
         default: C_AND = '0;
      endcase
   end
   //C_ANDI
   always_comb begin
      casez (data[31:0])
         32'b????????????????100?10????????01: C_ANDI = '1;
         default: C_ANDI = '0;
      endcase
   end
   //C_BEQZ
   always_comb begin
      casez (data[31:0])
         32'b????????????????110???????????01: C_BEQZ = '1;
         default: C_BEQZ = '0;
      endcase
   end
   //C_BNEZ
   always_comb begin
      casez (data[31:0])
         32'b????????????????111???????????01: C_BNEZ = '1;
         default: C_BNEZ = '0;
      endcase
   end
   //C_EBREAK
   always_comb begin
      casez (data[31:0])
         32'b????????????????1001000000000010: C_EBREAK = '1;
         default: C_EBREAK = '0;
      endcase
   end
   //C_J
   always_comb begin
      casez (data[31:0])
         32'b????????????????101???????????01: C_J = '1;
         default: C_J = '0;
      endcase
   end
   //C_JAL
   always_comb begin
      casez (data[31:0])
         32'b????????????????001???????????01: C_JAL = '1;
         default: C_JAL = '0;
      endcase
   end
   //C_JALR
   always_comb begin
      casez (data[31:0])
         32'b????????????????1001????10000010: C_JALR = '1;
         32'b????????????????10011????0000010: C_JALR = '1;
         32'b????????????????1001??1??0000010: C_JALR = '1;
         32'b????????????????1001???1?0000010: C_JALR = '1;
         32'b????????????????1001?1???0000010: C_JALR = '1;
         default: C_JALR = '0;
      endcase
   end
   //C_JR
   always_comb begin
      casez (data[31:0])
         32'b????????????????1000?????0000010: C_JR = '1;
         default: C_JR = '0;
      endcase
   end
   //C_LI
   always_comb begin
      casez (data[31:0])
         32'b????????????????010???????????01: C_LI = '1;
         default: C_LI = '0;
      endcase
   end
   //C_LUI
   always_comb begin
      casez (data[31:0])
         32'b????????????????011?1?????????01: C_LUI = '1;
         32'b????????????????011?????1?????01: C_LUI = '1;
         32'b????????????????011??1????????01: C_LUI = '1;
         32'b????????????????011????0??????01: C_LUI = '1;
         32'b????????????????011???1???????01: C_LUI = '1;
         default: C_LUI = '0;
      endcase
   end
   //C_LW
   always_comb begin
      casez (data[31:0])
         32'b????????????????010???????????00: C_LW = '1;
         default: C_LW = '0;
      endcase
   end
   //C_LWSP
   always_comb begin
      casez (data[31:0])
         32'b????????????????010????1??????10: C_LWSP = '1;
         32'b????????????????010???1???????10: C_LWSP = '1;
         32'b????????????????010??1????????10: C_LWSP = '1;
         32'b????????????????010?1?????????10: C_LWSP = '1;
         32'b????????????????010?????1?????10: C_LWSP = '1;
         default: C_LWSP = '0;
      endcase
   end
   //C_MV
   always_comb begin
      casez (data[31:0])
         32'b????????????????1000?????1????10: C_MV = '1;
         32'b????????????????1000???????1??10: C_MV = '1;
         32'b????????????????1000?????????110: C_MV = '1;
         32'b????????????????1000????????1?10: C_MV = '1;
         32'b????????????????1000??????1???10: C_MV = '1;
         default: C_MV = '0;
      endcase
   end
   //C_NOP
   always_comb begin
      casez (data[31:0])
         32'b????????????????000?00000?????01: C_NOP = '1;
         default: C_NOP = '0;
      endcase
   end
   //C_OR
   always_comb begin
      casez (data[31:0])
         32'b????????????????100011???10???01: C_OR = '1;
         default: C_OR = '0;
      endcase
   end
   //C_SUB
   always_comb begin
      casez (data[31:0])
         32'b????????????????100011???00???01: C_SUB = '1;
         default: C_SUB = '0;
      endcase
   end
   //C_SW
   always_comb begin
      casez (data[31:0])
         32'b????????????????110???????????00: C_SW = '1;
         default: C_SW = '0;
      endcase
   end
   //C_SWSP
   always_comb begin
      casez (data[31:0])
         32'b????????????????110???????????10: C_SWSP = '1;
         default: C_SWSP = '0;
      endcase
   end
   //C_XOR
   always_comb begin
      casez (data[31:0])
         32'b????????????????100011???01???01: C_XOR = '1;
         default: C_XOR = '0;
      endcase
   end
   //DIV
   always_comb begin
      casez (data[31:0])
         32'b0000001??????????100?????0110011: DIV = '1;
         default: DIV = '0;
      endcase
   end
   //DIVU
   always_comb begin
      casez (data[31:0])
         32'b0000001??????????101?????0110011: DIVU = '1;
         default: DIVU = '0;
      endcase
   end
   //EBREAK
   always_comb begin
      casez (data[31:0])
         32'b00000000000100000000000001110011: EBREAK = '1;
         default: EBREAK = '0;
      endcase
   end
   //ECALL
   always_comb begin
      casez (data[31:0])
         32'b00000000000000000000000001110011: ECALL = '1;
         default: ECALL = '0;
      endcase
   end
   //FENCE
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????0001111: FENCE = '1;
         default: FENCE = '0;
      endcase
   end
   //JAL
   always_comb begin
      casez (data[31:0])
         32'b?????????????????????????1101111: JAL = '1;
         default: JAL = '0;
      endcase
   end
   //JALR
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????1100111: JALR = '1;
         default: JALR = '0;
      endcase
   end
   //LB
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????0000011: LB = '1;
         default: LB = '0;
      endcase
   end
   //LBU
   always_comb begin
      casez (data[31:0])
         32'b?????????????????100?????0000011: LBU = '1;
         default: LBU = '0;
      endcase
   end
   //LH
   always_comb begin
      casez (data[31:0])
         32'b?????????????????001?????0000011: LH = '1;
         default: LH = '0;
      endcase
   end
   //LHU
   always_comb begin
      casez (data[31:0])
         32'b?????????????????101?????0000011: LHU = '1;
         default: LHU = '0;
      endcase
   end
   //LUI
   always_comb begin
      casez (data[31:0])
         32'b?????????????????????????0110111: LUI = '1;
         default: LUI = '0;
      endcase
   end
   //LW
   always_comb begin
      casez (data[31:0])
         32'b?????????????????010?????0000011: LW = '1;
         default: LW = '0;
      endcase
   end
   //MUL
   always_comb begin
      casez (data[31:0])
         32'b0000001??????????000?????0110011: MUL = '1;
         default: MUL = '0;
      endcase
   end
   //MULH
   always_comb begin
      casez (data[31:0])
         32'b0000001??????????001?????0110011: MULH = '1;
         default: MULH = '0;
      endcase
   end
   //MULHSU
   always_comb begin
      casez (data[31:0])
         32'b0000001??????????010?????0110011: MULHSU = '1;
         default: MULHSU = '0;
      endcase
   end
   //MULHU
   always_comb begin
      casez (data[31:0])
         32'b0000001??????????011?????0110011: MULHU = '1;
         default: MULHU = '0;
      endcase
   end
   //OR
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????110?????0110011: OR = '1;
         default: OR = '0;
      endcase
   end
   //ORI
   always_comb begin
      casez (data[31:0])
         32'b?????????????????110?????0010011: ORI = '1;
         default: ORI = '0;
      endcase
   end
   //REM
   always_comb begin
      casez (data[31:0])
         32'b0000001??????????110?????0110011: REM = '1;
         default: REM = '0;
      endcase
   end
   //REMU
   always_comb begin
      casez (data[31:0])
         32'b0000001??????????111?????0110011: REMU = '1;
         default: REMU = '0;
      endcase
   end
   //SB
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????0100011: SB = '1;
         default: SB = '0;
      endcase
   end
   //SH
   always_comb begin
      casez (data[31:0])
         32'b?????????????????001?????0100011: SH = '1;
         default: SH = '0;
      endcase
   end
   //SLL
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????001?????0110011: SLL = '1;
         default: SLL = '0;
      endcase
   end
   //SLT
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????010?????0110011: SLT = '1;
         default: SLT = '0;
      endcase
   end
   //SLTI
   always_comb begin
      casez (data[31:0])
         32'b?????????????????010?????0010011: SLTI = '1;
         default: SLTI = '0;
      endcase
   end
   //SLTIU
   always_comb begin
      casez (data[31:0])
         32'b?????????????????011?????0010011: SLTIU = '1;
         default: SLTIU = '0;
      endcase
   end
   //SLTU
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????011?????0110011: SLTU = '1;
         default: SLTU = '0;
      endcase
   end
   //SRA
   always_comb begin
      casez (data[31:0])
         32'b0100000??????????101?????0110011: SRA = '1;
         default: SRA = '0;
      endcase
   end
   //SRL
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????101?????0110011: SRL = '1;
         default: SRL = '0;
      endcase
   end
   //SUB
   always_comb begin
      casez (data[31:0])
         32'b0100000??????????000?????0110011: SUB = '1;
         default: SUB = '0;
      endcase
   end
   //SW
   always_comb begin
      casez (data[31:0])
         32'b?????????????????010?????0100011: SW = '1;
         default: SW = '0;
      endcase
   end
   //XOR
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????100?????0110011: XOR = '1;
         default: XOR = '0;
      endcase
   end
   //XORI
   always_comb begin
      casez (data[31:0])
         32'b?????????????????100?????0010011: XORI = '1;
         default: XORI = '0;
      endcase
   end
   //defined
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????000?????0110011: defined = '1;
         32'b?????????????????000?????0010011: defined = '1;
         32'b0000000??????????111?????0110011: defined = '1;
         32'b?????????????????111?????0010011: defined = '1;
         32'b?????????????????????????0010111: defined = '1;
         32'b?????????????????000?????1100011: defined = '1;
         32'b?????????????????101?????1100011: defined = '1;
         32'b?????????????????111?????1100011: defined = '1;
         32'b?????????????????100?????1100011: defined = '1;
         32'b?????????????????110?????1100011: defined = '1;
         32'b?????????????????001?????1100011: defined = '1;
         32'b????????????????1001????????1?10: defined = '1;
         32'b????????????????1001??????1???10: defined = '1;
         32'b????????????????1001???????1??10: defined = '1;
         32'b????????????????1001?????1????10: defined = '1;
         32'b????????????????1001?????????110: defined = '1;
         32'b????????????????000?1?????????01: defined = '1;
         32'b????????????????000??1????????01: defined = '1;
         32'b????????????????000?????1?????01: defined = '1;
         32'b????????????????000???1???????01: defined = '1;
         32'b????????????????000????1??????01: defined = '1;
         32'b????????????????011?00010?????01: defined = '1;
         32'b????????????????000???????????00: defined = '1;
         32'b????????????????100011???11???01: defined = '1;
         32'b????????????????100?10????????01: defined = '1;
         32'b????????????????110???????????01: defined = '1;
         32'b????????????????111???????????01: defined = '1;
         32'b????????????????1001000000000010: defined = '1;
         32'b????????????????101???????????01: defined = '1;
         32'b????????????????001???????????01: defined = '1;
         32'b????????????????1001????10000010: defined = '1;
         32'b????????????????10011????0000010: defined = '1;
         32'b????????????????1001??1??0000010: defined = '1;
         32'b????????????????1001???1?0000010: defined = '1;
         32'b????????????????1001?1???0000010: defined = '1;
         32'b????????????????1000?????0000010: defined = '1;
         32'b????????????????010???????????01: defined = '1;
         32'b????????????????011?1?????????01: defined = '1;
         32'b????????????????011?????1?????01: defined = '1;
         32'b????????????????011??1????????01: defined = '1;
         32'b????????????????011????0??????01: defined = '1;
         32'b????????????????011???1???????01: defined = '1;
         32'b????????????????010???????????00: defined = '1;
         32'b????????????????010????1??????10: defined = '1;
         32'b????????????????010???1???????10: defined = '1;
         32'b????????????????010??1????????10: defined = '1;
         32'b????????????????010?1?????????10: defined = '1;
         32'b????????????????010?????1?????10: defined = '1;
         32'b????????????????1000?????1????10: defined = '1;
         32'b????????????????1000???????1??10: defined = '1;
         32'b????????????????1000?????????110: defined = '1;
         32'b????????????????1000????????1?10: defined = '1;
         32'b????????????????1000??????1???10: defined = '1;
         32'b????????????????000?00000?????01: defined = '1;
         32'b????????????????100011???10???01: defined = '1;
         32'b????????????????100011???00???01: defined = '1;
         32'b????????????????110???????????00: defined = '1;
         32'b????????????????110???????????10: defined = '1;
         32'b????????????????100011???01???01: defined = '1;
         32'b0000001??????????100?????0110011: defined = '1;
         32'b0000001??????????101?????0110011: defined = '1;
         32'b00000000000100000000000001110011: defined = '1;
         32'b00000000000000000000000001110011: defined = '1;
         32'b?????????????????000?????0001111: defined = '1;
         32'b?????????????????????????1101111: defined = '1;
         32'b?????????????????000?????1100111: defined = '1;
         32'b?????????????????000?????0000011: defined = '1;
         32'b?????????????????100?????0000011: defined = '1;
         32'b?????????????????001?????0000011: defined = '1;
         32'b?????????????????101?????0000011: defined = '1;
         32'b?????????????????????????0110111: defined = '1;
         32'b?????????????????010?????0000011: defined = '1;
         32'b0000001??????????000?????0110011: defined = '1;
         32'b0000001??????????001?????0110011: defined = '1;
         32'b0000001??????????010?????0110011: defined = '1;
         32'b0000001??????????011?????0110011: defined = '1;
         32'b0000000??????????110?????0110011: defined = '1;
         32'b?????????????????110?????0010011: defined = '1;
         32'b0000001??????????110?????0110011: defined = '1;
         32'b0000001??????????111?????0110011: defined = '1;
         32'b?????????????????000?????0100011: defined = '1;
         32'b?????????????????001?????0100011: defined = '1;
         32'b0000000??????????001?????0110011: defined = '1;
         32'b0000000??????????010?????0110011: defined = '1;
         32'b?????????????????010?????0010011: defined = '1;
         32'b?????????????????011?????0010011: defined = '1;
         32'b0000000??????????011?????0110011: defined = '1;
         32'b0100000??????????101?????0110011: defined = '1;
         32'b0000000??????????101?????0110011: defined = '1;
         32'b0100000??????????000?????0110011: defined = '1;
         32'b?????????????????010?????0100011: defined = '1;
         32'b0000000??????????100?????0110011: defined = '1;
         32'b?????????????????100?????0010011: defined = '1;
         default: defined = '0;
      endcase
   end
   //compressed
   always_comb begin
      casez (data[31:0])
         32'b????????????????1001????????1?10: compressed = '1;
         32'b????????????????1001??????1???10: compressed = '1;
         32'b????????????????1001???????1??10: compressed = '1;
         32'b????????????????1001?????1????10: compressed = '1;
         32'b????????????????1001?????????110: compressed = '1;
         32'b????????????????000?1?????????01: compressed = '1;
         32'b????????????????000??1????????01: compressed = '1;
         32'b????????????????000?????1?????01: compressed = '1;
         32'b????????????????000???1???????01: compressed = '1;
         32'b????????????????000????1??????01: compressed = '1;
         32'b????????????????011?00010?????01: compressed = '1;
         32'b????????????????000???????????00: compressed = '1;
         32'b????????????????100011???11???01: compressed = '1;
         32'b????????????????100?10????????01: compressed = '1;
         32'b????????????????110???????????01: compressed = '1;
         32'b????????????????111???????????01: compressed = '1;
         32'b????????????????1001000000000010: compressed = '1;
         32'b????????????????101???????????01: compressed = '1;
         32'b????????????????001???????????01: compressed = '1;
         32'b????????????????1001????10000010: compressed = '1;
         32'b????????????????10011????0000010: compressed = '1;
         32'b????????????????1001??1??0000010: compressed = '1;
         32'b????????????????1001???1?0000010: compressed = '1;
         32'b????????????????1001?1???0000010: compressed = '1;
         32'b????????????????1000?????0000010: compressed = '1;
         32'b????????????????010???????????01: compressed = '1;
         32'b????????????????011?1?????????01: compressed = '1;
         32'b????????????????011?????1?????01: compressed = '1;
         32'b????????????????011??1????????01: compressed = '1;
         32'b????????????????011????0??????01: compressed = '1;
         32'b????????????????011???1???????01: compressed = '1;
         32'b????????????????010???????????00: compressed = '1;
         32'b????????????????010????1??????10: compressed = '1;
         32'b????????????????010???1???????10: compressed = '1;
         32'b????????????????010??1????????10: compressed = '1;
         32'b????????????????010?1?????????10: compressed = '1;
         32'b????????????????010?????1?????10: compressed = '1;
         32'b????????????????1000?????1????10: compressed = '1;
         32'b????????????????1000???????1??10: compressed = '1;
         32'b????????????????1000?????????110: compressed = '1;
         32'b????????????????1000????????1?10: compressed = '1;
         32'b????????????????1000??????1???10: compressed = '1;
         32'b????????????????000?00000?????01: compressed = '1;
         32'b????????????????100011???10???01: compressed = '1;
         32'b????????????????100011???00???01: compressed = '1;
         32'b????????????????110???????????00: compressed = '1;
         32'b????????????????110???????????10: compressed = '1;
         32'b????????????????100011???01???01: compressed = '1;
         default: compressed = '0;
      endcase
   end
   //bimm12hi
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????1100011: bimm12hi = '1;
         32'b?????????????????101?????1100011: bimm12hi = '1;
         32'b?????????????????111?????1100011: bimm12hi = '1;
         32'b?????????????????100?????1100011: bimm12hi = '1;
         32'b?????????????????110?????1100011: bimm12hi = '1;
         32'b?????????????????001?????1100011: bimm12hi = '1;
         default: bimm12hi = '0;
      endcase
   end
   //bimm12lo
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????1100011: bimm12lo = '1;
         32'b?????????????????101?????1100011: bimm12lo = '1;
         32'b?????????????????111?????1100011: bimm12lo = '1;
         32'b?????????????????100?????1100011: bimm12lo = '1;
         32'b?????????????????110?????1100011: bimm12lo = '1;
         32'b?????????????????001?????1100011: bimm12lo = '1;
         default: bimm12lo = '0;
      endcase
   end
   //c_bimm9hi
   always_comb begin
      casez (data[31:0])
         32'b????????????????110???????????01: c_bimm9hi = '1;
         32'b????????????????111???????????01: c_bimm9hi = '1;
         default: c_bimm9hi = '0;
      endcase
   end
   //c_bimm9lo
   always_comb begin
      casez (data[31:0])
         32'b????????????????110???????????01: c_bimm9lo = '1;
         32'b????????????????111???????????01: c_bimm9lo = '1;
         default: c_bimm9lo = '0;
      endcase
   end
   //c_imm12
   always_comb begin
      casez (data[31:0])
         32'b????????????????101???????????01: c_imm12 = '1;
         32'b????????????????001???????????01: c_imm12 = '1;
         default: c_imm12 = '0;
      endcase
   end
   //c_imm6hi
   always_comb begin
      casez (data[31:0])
         32'b????????????????100?10????????01: c_imm6hi = '1;
         32'b????????????????010???????????01: c_imm6hi = '1;
         default: c_imm6hi = '0;
      endcase
   end
   //c_imm6lo
   always_comb begin
      casez (data[31:0])
         32'b????????????????100?10????????01: c_imm6lo = '1;
         32'b????????????????010???????????01: c_imm6lo = '1;
         default: c_imm6lo = '0;
      endcase
   end
   //c_nzimm10hi
   always_comb begin
      casez (data[31:0])
         32'b????????????????011?00010?????01: c_nzimm10hi = '1;
         default: c_nzimm10hi = '0;
      endcase
   end
   //c_nzimm10lo
   always_comb begin
      casez (data[31:0])
         32'b????????????????011?00010?????01: c_nzimm10lo = '1;
         default: c_nzimm10lo = '0;
      endcase
   end
   //c_nzimm18hi
   always_comb begin
      casez (data[31:0])
         32'b????????????????011?1?????????01: c_nzimm18hi = '1;
         32'b????????????????011?????1?????01: c_nzimm18hi = '1;
         32'b????????????????011??1????????01: c_nzimm18hi = '1;
         32'b????????????????011????0??????01: c_nzimm18hi = '1;
         32'b????????????????011???1???????01: c_nzimm18hi = '1;
         32'b????????????????011?1?????????01: c_nzimm18hi = '1;
         32'b????????????????011?????1?????01: c_nzimm18hi = '1;
         32'b????????????????011??1????????01: c_nzimm18hi = '1;
         32'b????????????????011????0??????01: c_nzimm18hi = '1;
         32'b????????????????011???1???????01: c_nzimm18hi = '1;
         32'b????????????????011?1?????????01: c_nzimm18hi = '1;
         32'b????????????????011?????1?????01: c_nzimm18hi = '1;
         32'b????????????????011??1????????01: c_nzimm18hi = '1;
         32'b????????????????011????0??????01: c_nzimm18hi = '1;
         32'b????????????????011???1???????01: c_nzimm18hi = '1;
         32'b????????????????011?1?????????01: c_nzimm18hi = '1;
         32'b????????????????011?????1?????01: c_nzimm18hi = '1;
         32'b????????????????011??1????????01: c_nzimm18hi = '1;
         32'b????????????????011????0??????01: c_nzimm18hi = '1;
         32'b????????????????011???1???????01: c_nzimm18hi = '1;
         32'b????????????????011?1?????????01: c_nzimm18hi = '1;
         32'b????????????????011?????1?????01: c_nzimm18hi = '1;
         32'b????????????????011??1????????01: c_nzimm18hi = '1;
         32'b????????????????011????0??????01: c_nzimm18hi = '1;
         32'b????????????????011???1???????01: c_nzimm18hi = '1;
         default: c_nzimm18hi = '0;
      endcase
   end
   //c_nzimm18lo
   always_comb begin
      casez (data[31:0])
         32'b????????????????011?1?????????01: c_nzimm18lo = '1;
         32'b????????????????011?????1?????01: c_nzimm18lo = '1;
         32'b????????????????011??1????????01: c_nzimm18lo = '1;
         32'b????????????????011????0??????01: c_nzimm18lo = '1;
         32'b????????????????011???1???????01: c_nzimm18lo = '1;
         32'b????????????????011?1?????????01: c_nzimm18lo = '1;
         32'b????????????????011?????1?????01: c_nzimm18lo = '1;
         32'b????????????????011??1????????01: c_nzimm18lo = '1;
         32'b????????????????011????0??????01: c_nzimm18lo = '1;
         32'b????????????????011???1???????01: c_nzimm18lo = '1;
         32'b????????????????011?1?????????01: c_nzimm18lo = '1;
         32'b????????????????011?????1?????01: c_nzimm18lo = '1;
         32'b????????????????011??1????????01: c_nzimm18lo = '1;
         32'b????????????????011????0??????01: c_nzimm18lo = '1;
         32'b????????????????011???1???????01: c_nzimm18lo = '1;
         32'b????????????????011?1?????????01: c_nzimm18lo = '1;
         32'b????????????????011?????1?????01: c_nzimm18lo = '1;
         32'b????????????????011??1????????01: c_nzimm18lo = '1;
         32'b????????????????011????0??????01: c_nzimm18lo = '1;
         32'b????????????????011???1???????01: c_nzimm18lo = '1;
         32'b????????????????011?1?????????01: c_nzimm18lo = '1;
         32'b????????????????011?????1?????01: c_nzimm18lo = '1;
         32'b????????????????011??1????????01: c_nzimm18lo = '1;
         32'b????????????????011????0??????01: c_nzimm18lo = '1;
         32'b????????????????011???1???????01: c_nzimm18lo = '1;
         default: c_nzimm18lo = '0;
      endcase
   end
   //c_nzimm6hi
   always_comb begin
      casez (data[31:0])
         32'b????????????????000?1?????????01: c_nzimm6hi = '1;
         32'b????????????????000??1????????01: c_nzimm6hi = '1;
         32'b????????????????000?????1?????01: c_nzimm6hi = '1;
         32'b????????????????000???1???????01: c_nzimm6hi = '1;
         32'b????????????????000????1??????01: c_nzimm6hi = '1;
         32'b????????????????000?1?????????01: c_nzimm6hi = '1;
         32'b????????????????000??1????????01: c_nzimm6hi = '1;
         32'b????????????????000?????1?????01: c_nzimm6hi = '1;
         32'b????????????????000???1???????01: c_nzimm6hi = '1;
         32'b????????????????000????1??????01: c_nzimm6hi = '1;
         32'b????????????????000?1?????????01: c_nzimm6hi = '1;
         32'b????????????????000??1????????01: c_nzimm6hi = '1;
         32'b????????????????000?????1?????01: c_nzimm6hi = '1;
         32'b????????????????000???1???????01: c_nzimm6hi = '1;
         32'b????????????????000????1??????01: c_nzimm6hi = '1;
         32'b????????????????000?1?????????01: c_nzimm6hi = '1;
         32'b????????????????000??1????????01: c_nzimm6hi = '1;
         32'b????????????????000?????1?????01: c_nzimm6hi = '1;
         32'b????????????????000???1???????01: c_nzimm6hi = '1;
         32'b????????????????000????1??????01: c_nzimm6hi = '1;
         32'b????????????????000?1?????????01: c_nzimm6hi = '1;
         32'b????????????????000??1????????01: c_nzimm6hi = '1;
         32'b????????????????000?????1?????01: c_nzimm6hi = '1;
         32'b????????????????000???1???????01: c_nzimm6hi = '1;
         32'b????????????????000????1??????01: c_nzimm6hi = '1;
         32'b????????????????000?00000?????01: c_nzimm6hi = '1;
         default: c_nzimm6hi = '0;
      endcase
   end
   //c_nzimm6lo
   always_comb begin
      casez (data[31:0])
         32'b????????????????000?1?????????01: c_nzimm6lo = '1;
         32'b????????????????000??1????????01: c_nzimm6lo = '1;
         32'b????????????????000?????1?????01: c_nzimm6lo = '1;
         32'b????????????????000???1???????01: c_nzimm6lo = '1;
         32'b????????????????000????1??????01: c_nzimm6lo = '1;
         32'b????????????????000?1?????????01: c_nzimm6lo = '1;
         32'b????????????????000??1????????01: c_nzimm6lo = '1;
         32'b????????????????000?????1?????01: c_nzimm6lo = '1;
         32'b????????????????000???1???????01: c_nzimm6lo = '1;
         32'b????????????????000????1??????01: c_nzimm6lo = '1;
         32'b????????????????000?1?????????01: c_nzimm6lo = '1;
         32'b????????????????000??1????????01: c_nzimm6lo = '1;
         32'b????????????????000?????1?????01: c_nzimm6lo = '1;
         32'b????????????????000???1???????01: c_nzimm6lo = '1;
         32'b????????????????000????1??????01: c_nzimm6lo = '1;
         32'b????????????????000?1?????????01: c_nzimm6lo = '1;
         32'b????????????????000??1????????01: c_nzimm6lo = '1;
         32'b????????????????000?????1?????01: c_nzimm6lo = '1;
         32'b????????????????000???1???????01: c_nzimm6lo = '1;
         32'b????????????????000????1??????01: c_nzimm6lo = '1;
         32'b????????????????000?1?????????01: c_nzimm6lo = '1;
         32'b????????????????000??1????????01: c_nzimm6lo = '1;
         32'b????????????????000?????1?????01: c_nzimm6lo = '1;
         32'b????????????????000???1???????01: c_nzimm6lo = '1;
         32'b????????????????000????1??????01: c_nzimm6lo = '1;
         32'b????????????????000?00000?????01: c_nzimm6lo = '1;
         default: c_nzimm6lo = '0;
      endcase
   end
   //c_nzuimm10
   always_comb begin
      casez (data[31:0])
         32'b????????????????000???????????00: c_nzuimm10 = '1;
         default: c_nzuimm10 = '0;
      endcase
   end
   //c_rs2
   always_comb begin
      casez (data[31:0])
         32'b????????????????1001????????1?10: c_rs2 = '1;
         32'b????????????????1001??????1???10: c_rs2 = '1;
         32'b????????????????1001???????1??10: c_rs2 = '1;
         32'b????????????????1001?????1????10: c_rs2 = '1;
         32'b????????????????1001?????????110: c_rs2 = '1;
         32'b????????????????1001????????1?10: c_rs2 = '1;
         32'b????????????????1001??????1???10: c_rs2 = '1;
         32'b????????????????1001???????1??10: c_rs2 = '1;
         32'b????????????????1001?????1????10: c_rs2 = '1;
         32'b????????????????1001?????????110: c_rs2 = '1;
         32'b????????????????1001????????1?10: c_rs2 = '1;
         32'b????????????????1001??????1???10: c_rs2 = '1;
         32'b????????????????1001???????1??10: c_rs2 = '1;
         32'b????????????????1001?????1????10: c_rs2 = '1;
         32'b????????????????1001?????????110: c_rs2 = '1;
         32'b????????????????1001????????1?10: c_rs2 = '1;
         32'b????????????????1001??????1???10: c_rs2 = '1;
         32'b????????????????1001???????1??10: c_rs2 = '1;
         32'b????????????????1001?????1????10: c_rs2 = '1;
         32'b????????????????1001?????????110: c_rs2 = '1;
         32'b????????????????1001????????1?10: c_rs2 = '1;
         32'b????????????????1001??????1???10: c_rs2 = '1;
         32'b????????????????1001???????1??10: c_rs2 = '1;
         32'b????????????????1001?????1????10: c_rs2 = '1;
         32'b????????????????1001?????????110: c_rs2 = '1;
         32'b????????????????1000?????1????10: c_rs2 = '1;
         32'b????????????????1000???????1??10: c_rs2 = '1;
         32'b????????????????1000?????????110: c_rs2 = '1;
         32'b????????????????1000????????1?10: c_rs2 = '1;
         32'b????????????????1000??????1???10: c_rs2 = '1;
         32'b????????????????1000?????1????10: c_rs2 = '1;
         32'b????????????????1000???????1??10: c_rs2 = '1;
         32'b????????????????1000?????????110: c_rs2 = '1;
         32'b????????????????1000????????1?10: c_rs2 = '1;
         32'b????????????????1000??????1???10: c_rs2 = '1;
         32'b????????????????1000?????1????10: c_rs2 = '1;
         32'b????????????????1000???????1??10: c_rs2 = '1;
         32'b????????????????1000?????????110: c_rs2 = '1;
         32'b????????????????1000????????1?10: c_rs2 = '1;
         32'b????????????????1000??????1???10: c_rs2 = '1;
         32'b????????????????1000?????1????10: c_rs2 = '1;
         32'b????????????????1000???????1??10: c_rs2 = '1;
         32'b????????????????1000?????????110: c_rs2 = '1;
         32'b????????????????1000????????1?10: c_rs2 = '1;
         32'b????????????????1000??????1???10: c_rs2 = '1;
         32'b????????????????1000?????1????10: c_rs2 = '1;
         32'b????????????????1000???????1??10: c_rs2 = '1;
         32'b????????????????1000?????????110: c_rs2 = '1;
         32'b????????????????1000????????1?10: c_rs2 = '1;
         32'b????????????????1000??????1???10: c_rs2 = '1;
         32'b????????????????110???????????10: c_rs2 = '1;
         default: c_rs2 = '0;
      endcase
   end
   //c_uimm7hi
   always_comb begin
      casez (data[31:0])
         32'b????????????????010???????????00: c_uimm7hi = '1;
         32'b????????????????110???????????00: c_uimm7hi = '1;
         default: c_uimm7hi = '0;
      endcase
   end
   //c_uimm7lo
   always_comb begin
      casez (data[31:0])
         32'b????????????????010???????????00: c_uimm7lo = '1;
         32'b????????????????110???????????00: c_uimm7lo = '1;
         default: c_uimm7lo = '0;
      endcase
   end
   //c_uimm8sp_s
   always_comb begin
      casez (data[31:0])
         32'b????????????????110???????????10: c_uimm8sp_s = '1;
         default: c_uimm8sp_s = '0;
      endcase
   end
   //c_uimm8sphi
   always_comb begin
      casez (data[31:0])
         32'b????????????????010????1??????10: c_uimm8sphi = '1;
         32'b????????????????010???1???????10: c_uimm8sphi = '1;
         32'b????????????????010??1????????10: c_uimm8sphi = '1;
         32'b????????????????010?1?????????10: c_uimm8sphi = '1;
         32'b????????????????010?????1?????10: c_uimm8sphi = '1;
         32'b????????????????010????1??????10: c_uimm8sphi = '1;
         32'b????????????????010???1???????10: c_uimm8sphi = '1;
         32'b????????????????010??1????????10: c_uimm8sphi = '1;
         32'b????????????????010?1?????????10: c_uimm8sphi = '1;
         32'b????????????????010?????1?????10: c_uimm8sphi = '1;
         32'b????????????????010????1??????10: c_uimm8sphi = '1;
         32'b????????????????010???1???????10: c_uimm8sphi = '1;
         32'b????????????????010??1????????10: c_uimm8sphi = '1;
         32'b????????????????010?1?????????10: c_uimm8sphi = '1;
         32'b????????????????010?????1?????10: c_uimm8sphi = '1;
         32'b????????????????010????1??????10: c_uimm8sphi = '1;
         32'b????????????????010???1???????10: c_uimm8sphi = '1;
         32'b????????????????010??1????????10: c_uimm8sphi = '1;
         32'b????????????????010?1?????????10: c_uimm8sphi = '1;
         32'b????????????????010?????1?????10: c_uimm8sphi = '1;
         32'b????????????????010????1??????10: c_uimm8sphi = '1;
         32'b????????????????010???1???????10: c_uimm8sphi = '1;
         32'b????????????????010??1????????10: c_uimm8sphi = '1;
         32'b????????????????010?1?????????10: c_uimm8sphi = '1;
         32'b????????????????010?????1?????10: c_uimm8sphi = '1;
         default: c_uimm8sphi = '0;
      endcase
   end
   //c_uimm8splo
   always_comb begin
      casez (data[31:0])
         32'b????????????????010????1??????10: c_uimm8splo = '1;
         32'b????????????????010???1???????10: c_uimm8splo = '1;
         32'b????????????????010??1????????10: c_uimm8splo = '1;
         32'b????????????????010?1?????????10: c_uimm8splo = '1;
         32'b????????????????010?????1?????10: c_uimm8splo = '1;
         32'b????????????????010????1??????10: c_uimm8splo = '1;
         32'b????????????????010???1???????10: c_uimm8splo = '1;
         32'b????????????????010??1????????10: c_uimm8splo = '1;
         32'b????????????????010?1?????????10: c_uimm8splo = '1;
         32'b????????????????010?????1?????10: c_uimm8splo = '1;
         32'b????????????????010????1??????10: c_uimm8splo = '1;
         32'b????????????????010???1???????10: c_uimm8splo = '1;
         32'b????????????????010??1????????10: c_uimm8splo = '1;
         32'b????????????????010?1?????????10: c_uimm8splo = '1;
         32'b????????????????010?????1?????10: c_uimm8splo = '1;
         32'b????????????????010????1??????10: c_uimm8splo = '1;
         32'b????????????????010???1???????10: c_uimm8splo = '1;
         32'b????????????????010??1????????10: c_uimm8splo = '1;
         32'b????????????????010?1?????????10: c_uimm8splo = '1;
         32'b????????????????010?????1?????10: c_uimm8splo = '1;
         32'b????????????????010????1??????10: c_uimm8splo = '1;
         32'b????????????????010???1???????10: c_uimm8splo = '1;
         32'b????????????????010??1????????10: c_uimm8splo = '1;
         32'b????????????????010?1?????????10: c_uimm8splo = '1;
         32'b????????????????010?????1?????10: c_uimm8splo = '1;
         default: c_uimm8splo = '0;
      endcase
   end
   //fm
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????0001111: fm = '1;
         default: fm = '0;
      endcase
   end
   //imm12
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????0010011: imm12 = '1;
         32'b?????????????????111?????0010011: imm12 = '1;
         32'b?????????????????000?????1100111: imm12 = '1;
         32'b?????????????????000?????0000011: imm12 = '1;
         32'b?????????????????100?????0000011: imm12 = '1;
         32'b?????????????????001?????0000011: imm12 = '1;
         32'b?????????????????101?????0000011: imm12 = '1;
         32'b?????????????????010?????0000011: imm12 = '1;
         32'b?????????????????110?????0010011: imm12 = '1;
         32'b?????????????????010?????0010011: imm12 = '1;
         32'b?????????????????011?????0010011: imm12 = '1;
         32'b?????????????????100?????0010011: imm12 = '1;
         default: imm12 = '0;
      endcase
   end
   //imm12hi
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????0100011: imm12hi = '1;
         32'b?????????????????001?????0100011: imm12hi = '1;
         32'b?????????????????010?????0100011: imm12hi = '1;
         default: imm12hi = '0;
      endcase
   end
   //imm12lo
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????0100011: imm12lo = '1;
         32'b?????????????????001?????0100011: imm12lo = '1;
         32'b?????????????????010?????0100011: imm12lo = '1;
         default: imm12lo = '0;
      endcase
   end
   //imm20
   always_comb begin
      casez (data[31:0])
         32'b?????????????????????????0010111: imm20 = '1;
         32'b?????????????????????????0110111: imm20 = '1;
         default: imm20 = '0;
      endcase
   end
   //jimm20
   always_comb begin
      casez (data[31:0])
         32'b?????????????????????????1101111: jimm20 = '1;
         default: jimm20 = '0;
      endcase
   end
   //pred
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????0001111: pred = '1;
         default: pred = '0;
      endcase
   end
   //rd
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????000?????0110011: rd = '1;
         32'b?????????????????000?????0010011: rd = '1;
         32'b0000000??????????111?????0110011: rd = '1;
         32'b?????????????????111?????0010011: rd = '1;
         32'b?????????????????????????0010111: rd = '1;
         32'b????????????????010???????????01: rd = '1;
         32'b????????????????011?1?????????01: rd = '1;
         32'b????????????????011?????1?????01: rd = '1;
         32'b????????????????011??1????????01: rd = '1;
         32'b????????????????011????0??????01: rd = '1;
         32'b????????????????011???1???????01: rd = '1;
         32'b????????????????011?1?????????01: rd = '1;
         32'b????????????????011?????1?????01: rd = '1;
         32'b????????????????011??1????????01: rd = '1;
         32'b????????????????011????0??????01: rd = '1;
         32'b????????????????011???1???????01: rd = '1;
         32'b????????????????011?1?????????01: rd = '1;
         32'b????????????????011?????1?????01: rd = '1;
         32'b????????????????011??1????????01: rd = '1;
         32'b????????????????011????0??????01: rd = '1;
         32'b????????????????011???1???????01: rd = '1;
         32'b????????????????011?1?????????01: rd = '1;
         32'b????????????????011?????1?????01: rd = '1;
         32'b????????????????011??1????????01: rd = '1;
         32'b????????????????011????0??????01: rd = '1;
         32'b????????????????011???1???????01: rd = '1;
         32'b????????????????011?1?????????01: rd = '1;
         32'b????????????????011?????1?????01: rd = '1;
         32'b????????????????011??1????????01: rd = '1;
         32'b????????????????011????0??????01: rd = '1;
         32'b????????????????011???1???????01: rd = '1;
         32'b????????????????010????1??????10: rd = '1;
         32'b????????????????010???1???????10: rd = '1;
         32'b????????????????010??1????????10: rd = '1;
         32'b????????????????010?1?????????10: rd = '1;
         32'b????????????????010?????1?????10: rd = '1;
         32'b????????????????010????1??????10: rd = '1;
         32'b????????????????010???1???????10: rd = '1;
         32'b????????????????010??1????????10: rd = '1;
         32'b????????????????010?1?????????10: rd = '1;
         32'b????????????????010?????1?????10: rd = '1;
         32'b????????????????010????1??????10: rd = '1;
         32'b????????????????010???1???????10: rd = '1;
         32'b????????????????010??1????????10: rd = '1;
         32'b????????????????010?1?????????10: rd = '1;
         32'b????????????????010?????1?????10: rd = '1;
         32'b????????????????010????1??????10: rd = '1;
         32'b????????????????010???1???????10: rd = '1;
         32'b????????????????010??1????????10: rd = '1;
         32'b????????????????010?1?????????10: rd = '1;
         32'b????????????????010?????1?????10: rd = '1;
         32'b????????????????010????1??????10: rd = '1;
         32'b????????????????010???1???????10: rd = '1;
         32'b????????????????010??1????????10: rd = '1;
         32'b????????????????010?1?????????10: rd = '1;
         32'b????????????????010?????1?????10: rd = '1;
         32'b????????????????1000?????1????10: rd = '1;
         32'b????????????????1000???????1??10: rd = '1;
         32'b????????????????1000?????????110: rd = '1;
         32'b????????????????1000????????1?10: rd = '1;
         32'b????????????????1000??????1???10: rd = '1;
         32'b????????????????1000?????1????10: rd = '1;
         32'b????????????????1000???????1??10: rd = '1;
         32'b????????????????1000?????????110: rd = '1;
         32'b????????????????1000????????1?10: rd = '1;
         32'b????????????????1000??????1???10: rd = '1;
         32'b????????????????1000?????1????10: rd = '1;
         32'b????????????????1000???????1??10: rd = '1;
         32'b????????????????1000?????????110: rd = '1;
         32'b????????????????1000????????1?10: rd = '1;
         32'b????????????????1000??????1???10: rd = '1;
         32'b????????????????1000?????1????10: rd = '1;
         32'b????????????????1000???????1??10: rd = '1;
         32'b????????????????1000?????????110: rd = '1;
         32'b????????????????1000????????1?10: rd = '1;
         32'b????????????????1000??????1???10: rd = '1;
         32'b????????????????1000?????1????10: rd = '1;
         32'b????????????????1000???????1??10: rd = '1;
         32'b????????????????1000?????????110: rd = '1;
         32'b????????????????1000????????1?10: rd = '1;
         32'b????????????????1000??????1???10: rd = '1;
         32'b0000001??????????100?????0110011: rd = '1;
         32'b0000001??????????101?????0110011: rd = '1;
         32'b?????????????????000?????0001111: rd = '1;
         32'b?????????????????????????1101111: rd = '1;
         32'b?????????????????000?????1100111: rd = '1;
         32'b?????????????????000?????0000011: rd = '1;
         32'b?????????????????100?????0000011: rd = '1;
         32'b?????????????????001?????0000011: rd = '1;
         32'b?????????????????101?????0000011: rd = '1;
         32'b?????????????????????????0110111: rd = '1;
         32'b?????????????????010?????0000011: rd = '1;
         32'b0000001??????????000?????0110011: rd = '1;
         32'b0000001??????????001?????0110011: rd = '1;
         32'b0000001??????????010?????0110011: rd = '1;
         32'b0000001??????????011?????0110011: rd = '1;
         32'b0000000??????????110?????0110011: rd = '1;
         32'b?????????????????110?????0010011: rd = '1;
         32'b0000001??????????110?????0110011: rd = '1;
         32'b0000001??????????111?????0110011: rd = '1;
         32'b0000000??????????001?????0110011: rd = '1;
         32'b0000000??????????010?????0110011: rd = '1;
         32'b?????????????????010?????0010011: rd = '1;
         32'b?????????????????011?????0010011: rd = '1;
         32'b0000000??????????011?????0110011: rd = '1;
         32'b0100000??????????101?????0110011: rd = '1;
         32'b0000000??????????101?????0110011: rd = '1;
         32'b0100000??????????000?????0110011: rd = '1;
         32'b0000000??????????100?????0110011: rd = '1;
         32'b?????????????????100?????0010011: rd = '1;
         default: rd = '0;
      endcase
   end
   //rd_p
   always_comb begin
      casez (data[31:0])
         32'b????????????????000???????????00: rd_p = '1;
         32'b????????????????010???????????00: rd_p = '1;
         default: rd_p = '0;
      endcase
   end
   //rd_rs1
   always_comb begin
      casez (data[31:0])
         32'b????????????????1001????????1?10: rd_rs1 = '1;
         32'b????????????????1001??????1???10: rd_rs1 = '1;
         32'b????????????????1001???????1??10: rd_rs1 = '1;
         32'b????????????????1001?????1????10: rd_rs1 = '1;
         32'b????????????????1001?????????110: rd_rs1 = '1;
         32'b????????????????1001????????1?10: rd_rs1 = '1;
         32'b????????????????1001??????1???10: rd_rs1 = '1;
         32'b????????????????1001???????1??10: rd_rs1 = '1;
         32'b????????????????1001?????1????10: rd_rs1 = '1;
         32'b????????????????1001?????????110: rd_rs1 = '1;
         32'b????????????????1001????????1?10: rd_rs1 = '1;
         32'b????????????????1001??????1???10: rd_rs1 = '1;
         32'b????????????????1001???????1??10: rd_rs1 = '1;
         32'b????????????????1001?????1????10: rd_rs1 = '1;
         32'b????????????????1001?????????110: rd_rs1 = '1;
         32'b????????????????1001????????1?10: rd_rs1 = '1;
         32'b????????????????1001??????1???10: rd_rs1 = '1;
         32'b????????????????1001???????1??10: rd_rs1 = '1;
         32'b????????????????1001?????1????10: rd_rs1 = '1;
         32'b????????????????1001?????????110: rd_rs1 = '1;
         32'b????????????????1001????????1?10: rd_rs1 = '1;
         32'b????????????????1001??????1???10: rd_rs1 = '1;
         32'b????????????????1001???????1??10: rd_rs1 = '1;
         32'b????????????????1001?????1????10: rd_rs1 = '1;
         32'b????????????????1001?????????110: rd_rs1 = '1;
         32'b????????????????000?1?????????01: rd_rs1 = '1;
         32'b????????????????000??1????????01: rd_rs1 = '1;
         32'b????????????????000?????1?????01: rd_rs1 = '1;
         32'b????????????????000???1???????01: rd_rs1 = '1;
         32'b????????????????000????1??????01: rd_rs1 = '1;
         32'b????????????????000?1?????????01: rd_rs1 = '1;
         32'b????????????????000??1????????01: rd_rs1 = '1;
         32'b????????????????000?????1?????01: rd_rs1 = '1;
         32'b????????????????000???1???????01: rd_rs1 = '1;
         32'b????????????????000????1??????01: rd_rs1 = '1;
         32'b????????????????000?1?????????01: rd_rs1 = '1;
         32'b????????????????000??1????????01: rd_rs1 = '1;
         32'b????????????????000?????1?????01: rd_rs1 = '1;
         32'b????????????????000???1???????01: rd_rs1 = '1;
         32'b????????????????000????1??????01: rd_rs1 = '1;
         32'b????????????????000?1?????????01: rd_rs1 = '1;
         32'b????????????????000??1????????01: rd_rs1 = '1;
         32'b????????????????000?????1?????01: rd_rs1 = '1;
         32'b????????????????000???1???????01: rd_rs1 = '1;
         32'b????????????????000????1??????01: rd_rs1 = '1;
         32'b????????????????000?1?????????01: rd_rs1 = '1;
         32'b????????????????000??1????????01: rd_rs1 = '1;
         32'b????????????????000?????1?????01: rd_rs1 = '1;
         32'b????????????????000???1???????01: rd_rs1 = '1;
         32'b????????????????000????1??????01: rd_rs1 = '1;
         default: rd_rs1 = '0;
      endcase
   end
   //rd_rs1_p
   always_comb begin
      casez (data[31:0])
         32'b????????????????100011???11???01: rd_rs1_p = '1;
         32'b????????????????100?10????????01: rd_rs1_p = '1;
         32'b????????????????100011???10???01: rd_rs1_p = '1;
         32'b????????????????100011???00???01: rd_rs1_p = '1;
         32'b????????????????100011???01???01: rd_rs1_p = '1;
         default: rd_rs1_p = '0;
      endcase
   end
   //rs1
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????000?????0110011: rs1 = '1;
         32'b?????????????????000?????0010011: rs1 = '1;
         32'b0000000??????????111?????0110011: rs1 = '1;
         32'b?????????????????111?????0010011: rs1 = '1;
         32'b?????????????????000?????1100011: rs1 = '1;
         32'b?????????????????101?????1100011: rs1 = '1;
         32'b?????????????????111?????1100011: rs1 = '1;
         32'b?????????????????100?????1100011: rs1 = '1;
         32'b?????????????????110?????1100011: rs1 = '1;
         32'b?????????????????001?????1100011: rs1 = '1;
         32'b????????????????1000?????0000010: rs1 = '1;
         32'b0000001??????????100?????0110011: rs1 = '1;
         32'b0000001??????????101?????0110011: rs1 = '1;
         32'b?????????????????000?????0001111: rs1 = '1;
         32'b?????????????????000?????1100111: rs1 = '1;
         32'b?????????????????000?????0000011: rs1 = '1;
         32'b?????????????????100?????0000011: rs1 = '1;
         32'b?????????????????001?????0000011: rs1 = '1;
         32'b?????????????????101?????0000011: rs1 = '1;
         32'b?????????????????010?????0000011: rs1 = '1;
         32'b0000001??????????000?????0110011: rs1 = '1;
         32'b0000001??????????001?????0110011: rs1 = '1;
         32'b0000001??????????010?????0110011: rs1 = '1;
         32'b0000001??????????011?????0110011: rs1 = '1;
         32'b0000000??????????110?????0110011: rs1 = '1;
         32'b?????????????????110?????0010011: rs1 = '1;
         32'b0000001??????????110?????0110011: rs1 = '1;
         32'b0000001??????????111?????0110011: rs1 = '1;
         32'b?????????????????000?????0100011: rs1 = '1;
         32'b?????????????????001?????0100011: rs1 = '1;
         32'b0000000??????????001?????0110011: rs1 = '1;
         32'b0000000??????????010?????0110011: rs1 = '1;
         32'b?????????????????010?????0010011: rs1 = '1;
         32'b?????????????????011?????0010011: rs1 = '1;
         32'b0000000??????????011?????0110011: rs1 = '1;
         32'b0100000??????????101?????0110011: rs1 = '1;
         32'b0000000??????????101?????0110011: rs1 = '1;
         32'b0100000??????????000?????0110011: rs1 = '1;
         32'b?????????????????010?????0100011: rs1 = '1;
         32'b0000000??????????100?????0110011: rs1 = '1;
         32'b?????????????????100?????0010011: rs1 = '1;
         default: rs1 = '0;
      endcase
   end
   //rs1_p
   always_comb begin
      casez (data[31:0])
         32'b????????????????110???????????01: rs1_p = '1;
         32'b????????????????111???????????01: rs1_p = '1;
         32'b????????????????010???????????00: rs1_p = '1;
         32'b????????????????110???????????00: rs1_p = '1;
         default: rs1_p = '0;
      endcase
   end
   //rs2
   always_comb begin
      casez (data[31:0])
         32'b0000000??????????000?????0110011: rs2 = '1;
         32'b0000000??????????111?????0110011: rs2 = '1;
         32'b?????????????????000?????1100011: rs2 = '1;
         32'b?????????????????101?????1100011: rs2 = '1;
         32'b?????????????????111?????1100011: rs2 = '1;
         32'b?????????????????100?????1100011: rs2 = '1;
         32'b?????????????????110?????1100011: rs2 = '1;
         32'b?????????????????001?????1100011: rs2 = '1;
         32'b0000001??????????100?????0110011: rs2 = '1;
         32'b0000001??????????101?????0110011: rs2 = '1;
         32'b0000001??????????000?????0110011: rs2 = '1;
         32'b0000001??????????001?????0110011: rs2 = '1;
         32'b0000001??????????010?????0110011: rs2 = '1;
         32'b0000001??????????011?????0110011: rs2 = '1;
         32'b0000000??????????110?????0110011: rs2 = '1;
         32'b0000001??????????110?????0110011: rs2 = '1;
         32'b0000001??????????111?????0110011: rs2 = '1;
         32'b?????????????????000?????0100011: rs2 = '1;
         32'b?????????????????001?????0100011: rs2 = '1;
         32'b0000000??????????001?????0110011: rs2 = '1;
         32'b0000000??????????010?????0110011: rs2 = '1;
         32'b0000000??????????011?????0110011: rs2 = '1;
         32'b0100000??????????101?????0110011: rs2 = '1;
         32'b0000000??????????101?????0110011: rs2 = '1;
         32'b0100000??????????000?????0110011: rs2 = '1;
         32'b?????????????????010?????0100011: rs2 = '1;
         32'b0000000??????????100?????0110011: rs2 = '1;
         default: rs2 = '0;
      endcase
   end
   //rs2_p
   always_comb begin
      casez (data[31:0])
         32'b????????????????100011???11???01: rs2_p = '1;
         32'b????????????????100011???10???01: rs2_p = '1;
         32'b????????????????100011???00???01: rs2_p = '1;
         32'b????????????????110???????????00: rs2_p = '1;
         32'b????????????????100011???01???01: rs2_p = '1;
         default: rs2_p = '0;
      endcase
   end
   //succ
   always_comb begin
      casez (data[31:0])
         32'b?????????????????000?????0001111: succ = '1;
         default: succ = '0;
      endcase
   end
endmodule
