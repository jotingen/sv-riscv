function automatic logic riscv_decode_add(
input logic [31:0] data
);
logic ADD;
casez (data[31:0])
32'b0000000??????????000?????0110011: ADD = '1;
default: ADD = '0;
endcase
return ADD;
endfunction
function automatic logic riscv_decode_addi(
input logic [31:0] data
);
logic ADDI;
casez (data[31:0])
32'b?????????????????000?????0010011: ADDI = '1;
default: ADDI = '0;
endcase
return ADDI;
endfunction
function automatic logic riscv_decode_and(
input logic [31:0] data
);
logic AND;
casez (data[31:0])
32'b0000000??????????111?????0110011: AND = '1;
default: AND = '0;
endcase
return AND;
endfunction
function automatic logic riscv_decode_andi(
input logic [31:0] data
);
logic ANDI;
casez (data[31:0])
32'b?????????????????111?????0010011: ANDI = '1;
default: ANDI = '0;
endcase
return ANDI;
endfunction
function automatic logic riscv_decode_auipc(
input logic [31:0] data
);
logic AUIPC;
casez (data[31:0])
32'b?????????????????????????0010111: AUIPC = '1;
default: AUIPC = '0;
endcase
return AUIPC;
endfunction
function automatic logic riscv_decode_beq(
input logic [31:0] data
);
logic BEQ;
casez (data[31:0])
32'b?????????????????000?????1100011: BEQ = '1;
default: BEQ = '0;
endcase
return BEQ;
endfunction
function automatic logic riscv_decode_bge(
input logic [31:0] data
);
logic BGE;
casez (data[31:0])
32'b?????????????????101?????1100011: BGE = '1;
default: BGE = '0;
endcase
return BGE;
endfunction
function automatic logic riscv_decode_bgeu(
input logic [31:0] data
);
logic BGEU;
casez (data[31:0])
32'b?????????????????111?????1100011: BGEU = '1;
default: BGEU = '0;
endcase
return BGEU;
endfunction
function automatic logic riscv_decode_blt(
input logic [31:0] data
);
logic BLT;
casez (data[31:0])
32'b?????????????????100?????1100011: BLT = '1;
default: BLT = '0;
endcase
return BLT;
endfunction
function automatic logic riscv_decode_bltu(
input logic [31:0] data
);
logic BLTU;
casez (data[31:0])
32'b?????????????????110?????1100011: BLTU = '1;
default: BLTU = '0;
endcase
return BLTU;
endfunction
function automatic logic riscv_decode_bne(
input logic [31:0] data
);
logic BNE;
casez (data[31:0])
32'b?????????????????001?????1100011: BNE = '1;
default: BNE = '0;
endcase
return BNE;
endfunction
function automatic logic riscv_decode_c_add(
input logic [31:0] data
);
logic C_ADD;
casez (data[31:0])
32'b????????????????1001????????1?10: C_ADD = '1;
32'b????????????????1001??????1???10: C_ADD = '1;
32'b????????????????1001???????1??10: C_ADD = '1;
32'b????????????????1001?????1????10: C_ADD = '1;
32'b????????????????1001?????????110: C_ADD = '1;
default: C_ADD = '0;
endcase
return C_ADD;
endfunction
function automatic logic riscv_decode_c_addi(
input logic [31:0] data
);
logic C_ADDI;
casez (data[31:0])
32'b????????????????000?1?????????01: C_ADDI = '1;
32'b????????????????000??1????????01: C_ADDI = '1;
32'b????????????????000?????1?????01: C_ADDI = '1;
32'b????????????????000???1???????01: C_ADDI = '1;
32'b????????????????000????1??????01: C_ADDI = '1;
default: C_ADDI = '0;
endcase
return C_ADDI;
endfunction
function automatic logic riscv_decode_c_addi16sp(
input logic [31:0] data
);
logic C_ADDI16SP;
casez (data[31:0])
32'b????????????????011?00010?????01: C_ADDI16SP = '1;
default: C_ADDI16SP = '0;
endcase
return C_ADDI16SP;
endfunction
function automatic logic riscv_decode_c_addi4spn(
input logic [31:0] data
);
logic C_ADDI4SPN;
casez (data[31:0])
32'b????????????????000???????????00: C_ADDI4SPN = '1;
default: C_ADDI4SPN = '0;
endcase
return C_ADDI4SPN;
endfunction
function automatic logic riscv_decode_c_and(
input logic [31:0] data
);
logic C_AND;
casez (data[31:0])
32'b????????????????100011???11???01: C_AND = '1;
default: C_AND = '0;
endcase
return C_AND;
endfunction
function automatic logic riscv_decode_c_andi(
input logic [31:0] data
);
logic C_ANDI;
casez (data[31:0])
32'b????????????????100?10????????01: C_ANDI = '1;
default: C_ANDI = '0;
endcase
return C_ANDI;
endfunction
function automatic logic riscv_decode_c_beqz(
input logic [31:0] data
);
logic C_BEQZ;
casez (data[31:0])
32'b????????????????110???????????01: C_BEQZ = '1;
default: C_BEQZ = '0;
endcase
return C_BEQZ;
endfunction
function automatic logic riscv_decode_c_bnez(
input logic [31:0] data
);
logic C_BNEZ;
casez (data[31:0])
32'b????????????????111???????????01: C_BNEZ = '1;
default: C_BNEZ = '0;
endcase
return C_BNEZ;
endfunction
function automatic logic riscv_decode_c_ebreak(
input logic [31:0] data
);
logic C_EBREAK;
casez (data[31:0])
32'b????????????????1001000000000010: C_EBREAK = '1;
default: C_EBREAK = '0;
endcase
return C_EBREAK;
endfunction
function automatic logic riscv_decode_c_j(
input logic [31:0] data
);
logic C_J;
casez (data[31:0])
32'b????????????????101???????????01: C_J = '1;
default: C_J = '0;
endcase
return C_J;
endfunction
function automatic logic riscv_decode_c_jal(
input logic [31:0] data
);
logic C_JAL;
casez (data[31:0])
32'b????????????????001???????????01: C_JAL = '1;
default: C_JAL = '0;
endcase
return C_JAL;
endfunction
function automatic logic riscv_decode_c_jalr(
input logic [31:0] data
);
logic C_JALR;
casez (data[31:0])
32'b????????????????1001????10000010: C_JALR = '1;
32'b????????????????10011????0000010: C_JALR = '1;
32'b????????????????1001??1??0000010: C_JALR = '1;
32'b????????????????1001???1?0000010: C_JALR = '1;
32'b????????????????1001?1???0000010: C_JALR = '1;
default: C_JALR = '0;
endcase
return C_JALR;
endfunction
function automatic logic riscv_decode_c_jr(
input logic [31:0] data
);
logic C_JR;
casez (data[31:0])
32'b????????????????1000?????0000010: C_JR = '1;
default: C_JR = '0;
endcase
return C_JR;
endfunction
function automatic logic riscv_decode_c_li(
input logic [31:0] data
);
logic C_LI;
casez (data[31:0])
32'b????????????????010???????????01: C_LI = '1;
default: C_LI = '0;
endcase
return C_LI;
endfunction
function automatic logic riscv_decode_c_lui(
input logic [31:0] data
);
logic C_LUI;
casez (data[31:0])
32'b????????????????011?1?????????01: C_LUI = '1;
32'b????????????????011?????1?????01: C_LUI = '1;
32'b????????????????011??1????????01: C_LUI = '1;
32'b????????????????011????0??????01: C_LUI = '1;
32'b????????????????011???1???????01: C_LUI = '1;
default: C_LUI = '0;
endcase
return C_LUI;
endfunction
function automatic logic riscv_decode_c_lw(
input logic [31:0] data
);
logic C_LW;
casez (data[31:0])
32'b????????????????010???????????00: C_LW = '1;
default: C_LW = '0;
endcase
return C_LW;
endfunction
function automatic logic riscv_decode_c_lwsp(
input logic [31:0] data
);
logic C_LWSP;
casez (data[31:0])
32'b????????????????010????1??????10: C_LWSP = '1;
32'b????????????????010???1???????10: C_LWSP = '1;
32'b????????????????010??1????????10: C_LWSP = '1;
32'b????????????????010?1?????????10: C_LWSP = '1;
32'b????????????????010?????1?????10: C_LWSP = '1;
default: C_LWSP = '0;
endcase
return C_LWSP;
endfunction
function automatic logic riscv_decode_c_mv(
input logic [31:0] data
);
logic C_MV;
casez (data[31:0])
32'b????????????????1000?????1????10: C_MV = '1;
32'b????????????????1000???????1??10: C_MV = '1;
32'b????????????????1000?????????110: C_MV = '1;
32'b????????????????1000????????1?10: C_MV = '1;
32'b????????????????1000??????1???10: C_MV = '1;
default: C_MV = '0;
endcase
return C_MV;
endfunction
function automatic logic riscv_decode_c_nop(
input logic [31:0] data
);
logic C_NOP;
casez (data[31:0])
32'b????????????????000?00000?????01: C_NOP = '1;
default: C_NOP = '0;
endcase
return C_NOP;
endfunction
function automatic logic riscv_decode_c_or(
input logic [31:0] data
);
logic C_OR;
casez (data[31:0])
32'b????????????????100011???10???01: C_OR = '1;
default: C_OR = '0;
endcase
return C_OR;
endfunction
function automatic logic riscv_decode_c_slli(
input logic [31:0] data
);
logic C_SLLI;
casez (data[31:0])
32'b????????????????000???1???????10: C_SLLI = '1;
32'b????????????????000?????1?????10: C_SLLI = '1;
32'b????????????????000????1??????10: C_SLLI = '1;
32'b????????????????000?1?????????10: C_SLLI = '1;
32'b????????????????000??1????????10: C_SLLI = '1;
default: C_SLLI = '0;
endcase
return C_SLLI;
endfunction
function automatic logic riscv_decode_c_srai(
input logic [31:0] data
);
logic C_SRAI;
casez (data[31:0])
32'b????????????????100?01????????01: C_SRAI = '1;
default: C_SRAI = '0;
endcase
return C_SRAI;
endfunction
function automatic logic riscv_decode_c_srli(
input logic [31:0] data
);
logic C_SRLI;
casez (data[31:0])
32'b????????????????100?00????????01: C_SRLI = '1;
default: C_SRLI = '0;
endcase
return C_SRLI;
endfunction
function automatic logic riscv_decode_c_sub(
input logic [31:0] data
);
logic C_SUB;
casez (data[31:0])
32'b????????????????100011???00???01: C_SUB = '1;
default: C_SUB = '0;
endcase
return C_SUB;
endfunction
function automatic logic riscv_decode_c_sw(
input logic [31:0] data
);
logic C_SW;
casez (data[31:0])
32'b????????????????110???????????00: C_SW = '1;
default: C_SW = '0;
endcase
return C_SW;
endfunction
function automatic logic riscv_decode_c_swsp(
input logic [31:0] data
);
logic C_SWSP;
casez (data[31:0])
32'b????????????????110???????????10: C_SWSP = '1;
default: C_SWSP = '0;
endcase
return C_SWSP;
endfunction
function automatic logic riscv_decode_c_xor(
input logic [31:0] data
);
logic C_XOR;
casez (data[31:0])
32'b????????????????100011???01???01: C_XOR = '1;
default: C_XOR = '0;
endcase
return C_XOR;
endfunction
function automatic logic riscv_decode_div(
input logic [31:0] data
);
logic DIV;
casez (data[31:0])
32'b0000001??????????100?????0110011: DIV = '1;
default: DIV = '0;
endcase
return DIV;
endfunction
function automatic logic riscv_decode_divu(
input logic [31:0] data
);
logic DIVU;
casez (data[31:0])
32'b0000001??????????101?????0110011: DIVU = '1;
default: DIVU = '0;
endcase
return DIVU;
endfunction
function automatic logic riscv_decode_ebreak(
input logic [31:0] data
);
logic EBREAK;
casez (data[31:0])
32'b00000000000100000000000001110011: EBREAK = '1;
default: EBREAK = '0;
endcase
return EBREAK;
endfunction
function automatic logic riscv_decode_ecall(
input logic [31:0] data
);
logic ECALL;
casez (data[31:0])
32'b00000000000000000000000001110011: ECALL = '1;
default: ECALL = '0;
endcase
return ECALL;
endfunction
function automatic logic riscv_decode_fence(
input logic [31:0] data
);
logic FENCE;
casez (data[31:0])
32'b?????????????????000?????0001111: FENCE = '1;
default: FENCE = '0;
endcase
return FENCE;
endfunction
function automatic logic riscv_decode_jal(
input logic [31:0] data
);
logic JAL;
casez (data[31:0])
32'b?????????????????????????1101111: JAL = '1;
default: JAL = '0;
endcase
return JAL;
endfunction
function automatic logic riscv_decode_jalr(
input logic [31:0] data
);
logic JALR;
casez (data[31:0])
32'b?????????????????000?????1100111: JALR = '1;
default: JALR = '0;
endcase
return JALR;
endfunction
function automatic logic riscv_decode_lb(
input logic [31:0] data
);
logic LB;
casez (data[31:0])
32'b?????????????????000?????0000011: LB = '1;
default: LB = '0;
endcase
return LB;
endfunction
function automatic logic riscv_decode_lbu(
input logic [31:0] data
);
logic LBU;
casez (data[31:0])
32'b?????????????????100?????0000011: LBU = '1;
default: LBU = '0;
endcase
return LBU;
endfunction
function automatic logic riscv_decode_lh(
input logic [31:0] data
);
logic LH;
casez (data[31:0])
32'b?????????????????001?????0000011: LH = '1;
default: LH = '0;
endcase
return LH;
endfunction
function automatic logic riscv_decode_lhu(
input logic [31:0] data
);
logic LHU;
casez (data[31:0])
32'b?????????????????101?????0000011: LHU = '1;
default: LHU = '0;
endcase
return LHU;
endfunction
function automatic logic riscv_decode_lui(
input logic [31:0] data
);
logic LUI;
casez (data[31:0])
32'b?????????????????????????0110111: LUI = '1;
default: LUI = '0;
endcase
return LUI;
endfunction
function automatic logic riscv_decode_lw(
input logic [31:0] data
);
logic LW;
casez (data[31:0])
32'b?????????????????010?????0000011: LW = '1;
default: LW = '0;
endcase
return LW;
endfunction
function automatic logic riscv_decode_mul(
input logic [31:0] data
);
logic MUL;
casez (data[31:0])
32'b0000001??????????000?????0110011: MUL = '1;
default: MUL = '0;
endcase
return MUL;
endfunction
function automatic logic riscv_decode_mulh(
input logic [31:0] data
);
logic MULH;
casez (data[31:0])
32'b0000001??????????001?????0110011: MULH = '1;
default: MULH = '0;
endcase
return MULH;
endfunction
function automatic logic riscv_decode_mulhsu(
input logic [31:0] data
);
logic MULHSU;
casez (data[31:0])
32'b0000001??????????010?????0110011: MULHSU = '1;
default: MULHSU = '0;
endcase
return MULHSU;
endfunction
function automatic logic riscv_decode_mulhu(
input logic [31:0] data
);
logic MULHU;
casez (data[31:0])
32'b0000001??????????011?????0110011: MULHU = '1;
default: MULHU = '0;
endcase
return MULHU;
endfunction
function automatic logic riscv_decode_or(
input logic [31:0] data
);
logic OR;
casez (data[31:0])
32'b0000000??????????110?????0110011: OR = '1;
default: OR = '0;
endcase
return OR;
endfunction
function automatic logic riscv_decode_ori(
input logic [31:0] data
);
logic ORI;
casez (data[31:0])
32'b?????????????????110?????0010011: ORI = '1;
default: ORI = '0;
endcase
return ORI;
endfunction
function automatic logic riscv_decode_rem(
input logic [31:0] data
);
logic REM;
casez (data[31:0])
32'b0000001??????????110?????0110011: REM = '1;
default: REM = '0;
endcase
return REM;
endfunction
function automatic logic riscv_decode_remu(
input logic [31:0] data
);
logic REMU;
casez (data[31:0])
32'b0000001??????????111?????0110011: REMU = '1;
default: REMU = '0;
endcase
return REMU;
endfunction
function automatic logic riscv_decode_sb(
input logic [31:0] data
);
logic SB;
casez (data[31:0])
32'b?????????????????000?????0100011: SB = '1;
default: SB = '0;
endcase
return SB;
endfunction
function automatic logic riscv_decode_sh(
input logic [31:0] data
);
logic SH;
casez (data[31:0])
32'b?????????????????001?????0100011: SH = '1;
default: SH = '0;
endcase
return SH;
endfunction
function automatic logic riscv_decode_sll(
input logic [31:0] data
);
logic SLL;
casez (data[31:0])
32'b0000000??????????001?????0110011: SLL = '1;
default: SLL = '0;
endcase
return SLL;
endfunction
function automatic logic riscv_decode_slli(
input logic [31:0] data
);
logic SLLI;
casez (data[31:0])
32'b000000???????????001?????0010011: SLLI = '1;
default: SLLI = '0;
endcase
return SLLI;
endfunction
function automatic logic riscv_decode_slt(
input logic [31:0] data
);
logic SLT;
casez (data[31:0])
32'b0000000??????????010?????0110011: SLT = '1;
default: SLT = '0;
endcase
return SLT;
endfunction
function automatic logic riscv_decode_slti(
input logic [31:0] data
);
logic SLTI;
casez (data[31:0])
32'b?????????????????010?????0010011: SLTI = '1;
default: SLTI = '0;
endcase
return SLTI;
endfunction
function automatic logic riscv_decode_sltiu(
input logic [31:0] data
);
logic SLTIU;
casez (data[31:0])
32'b?????????????????011?????0010011: SLTIU = '1;
default: SLTIU = '0;
endcase
return SLTIU;
endfunction
function automatic logic riscv_decode_sltu(
input logic [31:0] data
);
logic SLTU;
casez (data[31:0])
32'b0000000??????????011?????0110011: SLTU = '1;
default: SLTU = '0;
endcase
return SLTU;
endfunction
function automatic logic riscv_decode_sra(
input logic [31:0] data
);
logic SRA;
casez (data[31:0])
32'b0100000??????????101?????0110011: SRA = '1;
default: SRA = '0;
endcase
return SRA;
endfunction
function automatic logic riscv_decode_srai(
input logic [31:0] data
);
logic SRAI;
casez (data[31:0])
32'b010000???????????101?????0010011: SRAI = '1;
default: SRAI = '0;
endcase
return SRAI;
endfunction
function automatic logic riscv_decode_srl(
input logic [31:0] data
);
logic SRL;
casez (data[31:0])
32'b0000000??????????101?????0110011: SRL = '1;
default: SRL = '0;
endcase
return SRL;
endfunction
function automatic logic riscv_decode_srli(
input logic [31:0] data
);
logic SRLI;
casez (data[31:0])
32'b000000???????????101?????0010011: SRLI = '1;
default: SRLI = '0;
endcase
return SRLI;
endfunction
function automatic logic riscv_decode_sub(
input logic [31:0] data
);
logic SUB;
casez (data[31:0])
32'b0100000??????????000?????0110011: SUB = '1;
default: SUB = '0;
endcase
return SUB;
endfunction
function automatic logic riscv_decode_sw(
input logic [31:0] data
);
logic SW;
casez (data[31:0])
32'b?????????????????010?????0100011: SW = '1;
default: SW = '0;
endcase
return SW;
endfunction
function automatic logic riscv_decode_xor(
input logic [31:0] data
);
logic XOR;
casez (data[31:0])
32'b0000000??????????100?????0110011: XOR = '1;
default: XOR = '0;
endcase
return XOR;
endfunction
function automatic logic riscv_decode_xori(
input logic [31:0] data
);
logic XORI;
casez (data[31:0])
32'b?????????????????100?????0010011: XORI = '1;
default: XORI = '0;
endcase
return XORI;
endfunction
function automatic logic [31:0] riscv_decode_add_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_addi_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_and_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_andi_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_auipc_mask(
);
return 32'h7f;
endfunction
function automatic logic [31:0] riscv_decode_beq_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_bge_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_bgeu_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_blt_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_bltu_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_bne_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_c_add_mask(
);
return 32'hf003;
endfunction
function automatic logic [31:0] riscv_decode_c_addi_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_addi16sp_mask(
);
return 32'hef83;
endfunction
function automatic logic [31:0] riscv_decode_c_addi4spn_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_and_mask(
);
return 32'hfc63;
endfunction
function automatic logic [31:0] riscv_decode_c_andi_mask(
);
return 32'hec03;
endfunction
function automatic logic [31:0] riscv_decode_c_beqz_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_bnez_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_ebreak_mask(
);
return 32'hffff;
endfunction
function automatic logic [31:0] riscv_decode_c_j_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_jal_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_jalr_mask(
);
return 32'hf07f;
endfunction
function automatic logic [31:0] riscv_decode_c_jr_mask(
);
return 32'hf07f;
endfunction
function automatic logic [31:0] riscv_decode_c_li_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_lui_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_lw_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_lwsp_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_mv_mask(
);
return 32'hf003;
endfunction
function automatic logic [31:0] riscv_decode_c_nop_mask(
);
return 32'hef83;
endfunction
function automatic logic [31:0] riscv_decode_c_or_mask(
);
return 32'hfc63;
endfunction
function automatic logic [31:0] riscv_decode_c_slli_mask(
);
return 32'hf003;
endfunction
function automatic logic [31:0] riscv_decode_c_srai_mask(
);
return 32'hfc03;
endfunction
function automatic logic [31:0] riscv_decode_c_srli_mask(
);
return 32'hfc03;
endfunction
function automatic logic [31:0] riscv_decode_c_sub_mask(
);
return 32'hfc63;
endfunction
function automatic logic [31:0] riscv_decode_c_sw_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_swsp_mask(
);
return 32'he003;
endfunction
function automatic logic [31:0] riscv_decode_c_xor_mask(
);
return 32'hfc63;
endfunction
function automatic logic [31:0] riscv_decode_div_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_divu_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_ebreak_mask(
);
return 32'hffffffff;
endfunction
function automatic logic [31:0] riscv_decode_ecall_mask(
);
return 32'hffffffff;
endfunction
function automatic logic [31:0] riscv_decode_fence_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_jal_mask(
);
return 32'h7f;
endfunction
function automatic logic [31:0] riscv_decode_jalr_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_lb_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_lbu_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_lh_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_lhu_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_lui_mask(
);
return 32'h7f;
endfunction
function automatic logic [31:0] riscv_decode_lw_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_mul_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_mulh_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_mulhsu_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_mulhu_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_or_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_ori_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_rem_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_remu_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_sb_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_sh_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_sll_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_slli_mask(
);
return 32'hfc00707f;
endfunction
function automatic logic [31:0] riscv_decode_slt_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_slti_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_sltiu_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_sltu_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_sra_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_srai_mask(
);
return 32'hfc00707f;
endfunction
function automatic logic [31:0] riscv_decode_srl_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_srli_mask(
);
return 32'hfc00707f;
endfunction
function automatic logic [31:0] riscv_decode_sub_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_sw_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_xor_mask(
);
return 32'hfe00707f;
endfunction
function automatic logic [31:0] riscv_decode_xori_mask(
);
return 32'h707f;
endfunction
function automatic logic [31:0] riscv_decode_add_match(
);
return 32'h33;
endfunction
function automatic logic [31:0] riscv_decode_addi_match(
);
return 32'h13;
endfunction
function automatic logic [31:0] riscv_decode_and_match(
);
return 32'h7033;
endfunction
function automatic logic [31:0] riscv_decode_andi_match(
);
return 32'h7013;
endfunction
function automatic logic [31:0] riscv_decode_auipc_match(
);
return 32'h17;
endfunction
function automatic logic [31:0] riscv_decode_beq_match(
);
return 32'h63;
endfunction
function automatic logic [31:0] riscv_decode_bge_match(
);
return 32'h5063;
endfunction
function automatic logic [31:0] riscv_decode_bgeu_match(
);
return 32'h7063;
endfunction
function automatic logic [31:0] riscv_decode_blt_match(
);
return 32'h4063;
endfunction
function automatic logic [31:0] riscv_decode_bltu_match(
);
return 32'h6063;
endfunction
function automatic logic [31:0] riscv_decode_bne_match(
);
return 32'h1063;
endfunction
function automatic logic [31:0] riscv_decode_c_add_match(
);
return 32'h9002;
endfunction
function automatic logic [31:0] riscv_decode_c_addi_match(
);
return 32'h1;
endfunction
function automatic logic [31:0] riscv_decode_c_addi16sp_match(
);
return 32'h6101;
endfunction
function automatic logic [31:0] riscv_decode_c_addi4spn_match(
);
return 32'h0;
endfunction
function automatic logic [31:0] riscv_decode_c_and_match(
);
return 32'h8c61;
endfunction
function automatic logic [31:0] riscv_decode_c_andi_match(
);
return 32'h8801;
endfunction
function automatic logic [31:0] riscv_decode_c_beqz_match(
);
return 32'hc001;
endfunction
function automatic logic [31:0] riscv_decode_c_bnez_match(
);
return 32'he001;
endfunction
function automatic logic [31:0] riscv_decode_c_ebreak_match(
);
return 32'h9002;
endfunction
function automatic logic [31:0] riscv_decode_c_j_match(
);
return 32'ha001;
endfunction
function automatic logic [31:0] riscv_decode_c_jal_match(
);
return 32'h2001;
endfunction
function automatic logic [31:0] riscv_decode_c_jalr_match(
);
return 32'h9002;
endfunction
function automatic logic [31:0] riscv_decode_c_jr_match(
);
return 32'h8002;
endfunction
function automatic logic [31:0] riscv_decode_c_li_match(
);
return 32'h4001;
endfunction
function automatic logic [31:0] riscv_decode_c_lui_match(
);
return 32'h6001;
endfunction
function automatic logic [31:0] riscv_decode_c_lw_match(
);
return 32'h4000;
endfunction
function automatic logic [31:0] riscv_decode_c_lwsp_match(
);
return 32'h4002;
endfunction
function automatic logic [31:0] riscv_decode_c_mv_match(
);
return 32'h8002;
endfunction
function automatic logic [31:0] riscv_decode_c_nop_match(
);
return 32'h1;
endfunction
function automatic logic [31:0] riscv_decode_c_or_match(
);
return 32'h8c41;
endfunction
function automatic logic [31:0] riscv_decode_c_slli_match(
);
return 32'h2;
endfunction
function automatic logic [31:0] riscv_decode_c_srai_match(
);
return 32'h8401;
endfunction
function automatic logic [31:0] riscv_decode_c_srli_match(
);
return 32'h8001;
endfunction
function automatic logic [31:0] riscv_decode_c_sub_match(
);
return 32'h8c01;
endfunction
function automatic logic [31:0] riscv_decode_c_sw_match(
);
return 32'hc000;
endfunction
function automatic logic [31:0] riscv_decode_c_swsp_match(
);
return 32'hc002;
endfunction
function automatic logic [31:0] riscv_decode_c_xor_match(
);
return 32'h8c21;
endfunction
function automatic logic [31:0] riscv_decode_div_match(
);
return 32'h2004033;
endfunction
function automatic logic [31:0] riscv_decode_divu_match(
);
return 32'h2005033;
endfunction
function automatic logic [31:0] riscv_decode_ebreak_match(
);
return 32'h100073;
endfunction
function automatic logic [31:0] riscv_decode_ecall_match(
);
return 32'h73;
endfunction
function automatic logic [31:0] riscv_decode_fence_match(
);
return 32'hf;
endfunction
function automatic logic [31:0] riscv_decode_jal_match(
);
return 32'h6f;
endfunction
function automatic logic [31:0] riscv_decode_jalr_match(
);
return 32'h67;
endfunction
function automatic logic [31:0] riscv_decode_lb_match(
);
return 32'h3;
endfunction
function automatic logic [31:0] riscv_decode_lbu_match(
);
return 32'h4003;
endfunction
function automatic logic [31:0] riscv_decode_lh_match(
);
return 32'h1003;
endfunction
function automatic logic [31:0] riscv_decode_lhu_match(
);
return 32'h5003;
endfunction
function automatic logic [31:0] riscv_decode_lui_match(
);
return 32'h37;
endfunction
function automatic logic [31:0] riscv_decode_lw_match(
);
return 32'h2003;
endfunction
function automatic logic [31:0] riscv_decode_mul_match(
);
return 32'h2000033;
endfunction
function automatic logic [31:0] riscv_decode_mulh_match(
);
return 32'h2001033;
endfunction
function automatic logic [31:0] riscv_decode_mulhsu_match(
);
return 32'h2002033;
endfunction
function automatic logic [31:0] riscv_decode_mulhu_match(
);
return 32'h2003033;
endfunction
function automatic logic [31:0] riscv_decode_or_match(
);
return 32'h6033;
endfunction
function automatic logic [31:0] riscv_decode_ori_match(
);
return 32'h6013;
endfunction
function automatic logic [31:0] riscv_decode_rem_match(
);
return 32'h2006033;
endfunction
function automatic logic [31:0] riscv_decode_remu_match(
);
return 32'h2007033;
endfunction
function automatic logic [31:0] riscv_decode_sb_match(
);
return 32'h23;
endfunction
function automatic logic [31:0] riscv_decode_sh_match(
);
return 32'h1023;
endfunction
function automatic logic [31:0] riscv_decode_sll_match(
);
return 32'h1033;
endfunction
function automatic logic [31:0] riscv_decode_slli_match(
);
return 32'h1013;
endfunction
function automatic logic [31:0] riscv_decode_slt_match(
);
return 32'h2033;
endfunction
function automatic logic [31:0] riscv_decode_slti_match(
);
return 32'h2013;
endfunction
function automatic logic [31:0] riscv_decode_sltiu_match(
);
return 32'h3013;
endfunction
function automatic logic [31:0] riscv_decode_sltu_match(
);
return 32'h3033;
endfunction
function automatic logic [31:0] riscv_decode_sra_match(
);
return 32'h40005033;
endfunction
function automatic logic [31:0] riscv_decode_srai_match(
);
return 32'h40005013;
endfunction
function automatic logic [31:0] riscv_decode_srl_match(
);
return 32'h5033;
endfunction
function automatic logic [31:0] riscv_decode_srli_match(
);
return 32'h5013;
endfunction
function automatic logic [31:0] riscv_decode_sub_match(
);
return 32'h40000033;
endfunction
function automatic logic [31:0] riscv_decode_sw_match(
);
return 32'h2023;
endfunction
function automatic logic [31:0] riscv_decode_xor_match(
);
return 32'h4033;
endfunction
function automatic logic [31:0] riscv_decode_xori_match(
);
return 32'h4013;
endfunction
function automatic logic riscv_decode_defined(
input logic [31:0] data
);
logic defined;
casez (data[31:0])
32'b0000000??????????000?????0110011: defined = '1;
32'b?????????????????000?????0010011: defined = '1;
32'b0000000??????????111?????0110011: defined = '1;
32'b?????????????????111?????0010011: defined = '1;
32'b?????????????????????????0010111: defined = '1;
32'b?????????????????000?????1100011: defined = '1;
32'b?????????????????101?????1100011: defined = '1;
32'b?????????????????111?????1100011: defined = '1;
32'b?????????????????100?????1100011: defined = '1;
32'b?????????????????110?????1100011: defined = '1;
32'b?????????????????001?????1100011: defined = '1;
32'b????????????????1001????????1?10: defined = '1;
32'b????????????????1001??????1???10: defined = '1;
32'b????????????????1001???????1??10: defined = '1;
32'b????????????????1001?????1????10: defined = '1;
32'b????????????????1001?????????110: defined = '1;
32'b????????????????000?1?????????01: defined = '1;
32'b????????????????000??1????????01: defined = '1;
32'b????????????????000?????1?????01: defined = '1;
32'b????????????????000???1???????01: defined = '1;
32'b????????????????000????1??????01: defined = '1;
32'b????????????????011?00010?????01: defined = '1;
32'b????????????????000???????????00: defined = '1;
32'b????????????????100011???11???01: defined = '1;
32'b????????????????100?10????????01: defined = '1;
32'b????????????????110???????????01: defined = '1;
32'b????????????????111???????????01: defined = '1;
32'b????????????????1001000000000010: defined = '1;
32'b????????????????101???????????01: defined = '1;
32'b????????????????001???????????01: defined = '1;
32'b????????????????1001????10000010: defined = '1;
32'b????????????????10011????0000010: defined = '1;
32'b????????????????1001??1??0000010: defined = '1;
32'b????????????????1001???1?0000010: defined = '1;
32'b????????????????1001?1???0000010: defined = '1;
32'b????????????????1000?????0000010: defined = '1;
32'b????????????????010???????????01: defined = '1;
32'b????????????????011?1?????????01: defined = '1;
32'b????????????????011?????1?????01: defined = '1;
32'b????????????????011??1????????01: defined = '1;
32'b????????????????011????0??????01: defined = '1;
32'b????????????????011???1???????01: defined = '1;
32'b????????????????010???????????00: defined = '1;
32'b????????????????010????1??????10: defined = '1;
32'b????????????????010???1???????10: defined = '1;
32'b????????????????010??1????????10: defined = '1;
32'b????????????????010?1?????????10: defined = '1;
32'b????????????????010?????1?????10: defined = '1;
32'b????????????????1000?????1????10: defined = '1;
32'b????????????????1000???????1??10: defined = '1;
32'b????????????????1000?????????110: defined = '1;
32'b????????????????1000????????1?10: defined = '1;
32'b????????????????1000??????1???10: defined = '1;
32'b????????????????000?00000?????01: defined = '1;
32'b????????????????100011???10???01: defined = '1;
32'b????????????????000???1???????10: defined = '1;
32'b????????????????000?????1?????10: defined = '1;
32'b????????????????000????1??????10: defined = '1;
32'b????????????????000?1?????????10: defined = '1;
32'b????????????????000??1????????10: defined = '1;
32'b????????????????100?01????????01: defined = '1;
32'b????????????????100?00????????01: defined = '1;
32'b????????????????100011???00???01: defined = '1;
32'b????????????????110???????????00: defined = '1;
32'b????????????????110???????????10: defined = '1;
32'b????????????????100011???01???01: defined = '1;
32'b0000001??????????100?????0110011: defined = '1;
32'b0000001??????????101?????0110011: defined = '1;
32'b00000000000100000000000001110011: defined = '1;
32'b00000000000000000000000001110011: defined = '1;
32'b?????????????????000?????0001111: defined = '1;
32'b?????????????????????????1101111: defined = '1;
32'b?????????????????000?????1100111: defined = '1;
32'b?????????????????000?????0000011: defined = '1;
32'b?????????????????100?????0000011: defined = '1;
32'b?????????????????001?????0000011: defined = '1;
32'b?????????????????101?????0000011: defined = '1;
32'b?????????????????????????0110111: defined = '1;
32'b?????????????????010?????0000011: defined = '1;
32'b0000001??????????000?????0110011: defined = '1;
32'b0000001??????????001?????0110011: defined = '1;
32'b0000001??????????010?????0110011: defined = '1;
32'b0000001??????????011?????0110011: defined = '1;
32'b0000000??????????110?????0110011: defined = '1;
32'b?????????????????110?????0010011: defined = '1;
32'b0000001??????????110?????0110011: defined = '1;
32'b0000001??????????111?????0110011: defined = '1;
32'b?????????????????000?????0100011: defined = '1;
32'b?????????????????001?????0100011: defined = '1;
32'b0000000??????????001?????0110011: defined = '1;
32'b000000???????????001?????0010011: defined = '1;
32'b0000000??????????010?????0110011: defined = '1;
32'b?????????????????010?????0010011: defined = '1;
32'b?????????????????011?????0010011: defined = '1;
32'b0000000??????????011?????0110011: defined = '1;
32'b0100000??????????101?????0110011: defined = '1;
32'b010000???????????101?????0010011: defined = '1;
32'b0000000??????????101?????0110011: defined = '1;
32'b000000???????????101?????0010011: defined = '1;
32'b0100000??????????000?????0110011: defined = '1;
32'b?????????????????010?????0100011: defined = '1;
32'b0000000??????????100?????0110011: defined = '1;
32'b?????????????????100?????0010011: defined = '1;
default: defined = '0;
endcase
return defined;
endfunction
function automatic logic riscv_decode_compressed(
input logic [31:0] data
);
logic compressed;
casez (data[31:0])
32'b????????????????1001????????1?10: compressed = '1;
32'b????????????????1001??????1???10: compressed = '1;
32'b????????????????1001???????1??10: compressed = '1;
32'b????????????????1001?????1????10: compressed = '1;
32'b????????????????1001?????????110: compressed = '1;
32'b????????????????000?1?????????01: compressed = '1;
32'b????????????????000??1????????01: compressed = '1;
32'b????????????????000?????1?????01: compressed = '1;
32'b????????????????000???1???????01: compressed = '1;
32'b????????????????000????1??????01: compressed = '1;
32'b????????????????011?00010?????01: compressed = '1;
32'b????????????????000???????????00: compressed = '1;
32'b????????????????100011???11???01: compressed = '1;
32'b????????????????100?10????????01: compressed = '1;
32'b????????????????110???????????01: compressed = '1;
32'b????????????????111???????????01: compressed = '1;
32'b????????????????1001000000000010: compressed = '1;
32'b????????????????101???????????01: compressed = '1;
32'b????????????????001???????????01: compressed = '1;
32'b????????????????1001????10000010: compressed = '1;
32'b????????????????10011????0000010: compressed = '1;
32'b????????????????1001??1??0000010: compressed = '1;
32'b????????????????1001???1?0000010: compressed = '1;
32'b????????????????1001?1???0000010: compressed = '1;
32'b????????????????1000?????0000010: compressed = '1;
32'b????????????????010???????????01: compressed = '1;
32'b????????????????011?1?????????01: compressed = '1;
32'b????????????????011?????1?????01: compressed = '1;
32'b????????????????011??1????????01: compressed = '1;
32'b????????????????011????0??????01: compressed = '1;
32'b????????????????011???1???????01: compressed = '1;
32'b????????????????010???????????00: compressed = '1;
32'b????????????????010????1??????10: compressed = '1;
32'b????????????????010???1???????10: compressed = '1;
32'b????????????????010??1????????10: compressed = '1;
32'b????????????????010?1?????????10: compressed = '1;
32'b????????????????010?????1?????10: compressed = '1;
32'b????????????????1000?????1????10: compressed = '1;
32'b????????????????1000???????1??10: compressed = '1;
32'b????????????????1000?????????110: compressed = '1;
32'b????????????????1000????????1?10: compressed = '1;
32'b????????????????1000??????1???10: compressed = '1;
32'b????????????????000?00000?????01: compressed = '1;
32'b????????????????100011???10???01: compressed = '1;
32'b????????????????000???1???????10: compressed = '1;
32'b????????????????000?????1?????10: compressed = '1;
32'b????????????????000????1??????10: compressed = '1;
32'b????????????????000?1?????????10: compressed = '1;
32'b????????????????000??1????????10: compressed = '1;
32'b????????????????100?01????????01: compressed = '1;
32'b????????????????100?00????????01: compressed = '1;
32'b????????????????100011???00???01: compressed = '1;
32'b????????????????110???????????00: compressed = '1;
32'b????????????????110???????????10: compressed = '1;
32'b????????????????100011???01???01: compressed = '1;
default: compressed = '0;
endcase
return compressed;
endfunction
function automatic logic riscv_decode_bimm12hi(
input logic [31:0] data
);
logic bimm12hi;
casez (data[31:0])
32'b?????????????????000?????1100011: bimm12hi = '1;
32'b?????????????????101?????1100011: bimm12hi = '1;
32'b?????????????????111?????1100011: bimm12hi = '1;
32'b?????????????????100?????1100011: bimm12hi = '1;
32'b?????????????????110?????1100011: bimm12hi = '1;
32'b?????????????????001?????1100011: bimm12hi = '1;
default: bimm12hi = '0;
endcase
return bimm12hi;
endfunction
function automatic logic riscv_decode_bimm12lo(
input logic [31:0] data
);
logic bimm12lo;
casez (data[31:0])
32'b?????????????????000?????1100011: bimm12lo = '1;
32'b?????????????????101?????1100011: bimm12lo = '1;
32'b?????????????????111?????1100011: bimm12lo = '1;
32'b?????????????????100?????1100011: bimm12lo = '1;
32'b?????????????????110?????1100011: bimm12lo = '1;
32'b?????????????????001?????1100011: bimm12lo = '1;
default: bimm12lo = '0;
endcase
return bimm12lo;
endfunction
function automatic logic riscv_decode_c_bimm9hi(
input logic [31:0] data
);
logic c_bimm9hi;
casez (data[31:0])
32'b????????????????110???????????01: c_bimm9hi = '1;
32'b????????????????111???????????01: c_bimm9hi = '1;
default: c_bimm9hi = '0;
endcase
return c_bimm9hi;
endfunction
function automatic logic riscv_decode_c_bimm9lo(
input logic [31:0] data
);
logic c_bimm9lo;
casez (data[31:0])
32'b????????????????110???????????01: c_bimm9lo = '1;
32'b????????????????111???????????01: c_bimm9lo = '1;
default: c_bimm9lo = '0;
endcase
return c_bimm9lo;
endfunction
function automatic logic riscv_decode_c_imm12(
input logic [31:0] data
);
logic c_imm12;
casez (data[31:0])
32'b????????????????101???????????01: c_imm12 = '1;
32'b????????????????001???????????01: c_imm12 = '1;
default: c_imm12 = '0;
endcase
return c_imm12;
endfunction
function automatic logic riscv_decode_c_imm6hi(
input logic [31:0] data
);
logic c_imm6hi;
casez (data[31:0])
32'b????????????????100?10????????01: c_imm6hi = '1;
32'b????????????????010???????????01: c_imm6hi = '1;
default: c_imm6hi = '0;
endcase
return c_imm6hi;
endfunction
function automatic logic riscv_decode_c_imm6lo(
input logic [31:0] data
);
logic c_imm6lo;
casez (data[31:0])
32'b????????????????100?10????????01: c_imm6lo = '1;
32'b????????????????010???????????01: c_imm6lo = '1;
default: c_imm6lo = '0;
endcase
return c_imm6lo;
endfunction
function automatic logic riscv_decode_c_nzimm10hi(
input logic [31:0] data
);
logic c_nzimm10hi;
casez (data[31:0])
32'b????????????????011?00010?????01: c_nzimm10hi = '1;
default: c_nzimm10hi = '0;
endcase
return c_nzimm10hi;
endfunction
function automatic logic riscv_decode_c_nzimm10lo(
input logic [31:0] data
);
logic c_nzimm10lo;
casez (data[31:0])
32'b????????????????011?00010?????01: c_nzimm10lo = '1;
default: c_nzimm10lo = '0;
endcase
return c_nzimm10lo;
endfunction
function automatic logic riscv_decode_c_nzimm18hi(
input logic [31:0] data
);
logic c_nzimm18hi;
casez (data[31:0])
32'b????????????????011?1?????????01: c_nzimm18hi = '1;
32'b????????????????011?????1?????01: c_nzimm18hi = '1;
32'b????????????????011??1????????01: c_nzimm18hi = '1;
32'b????????????????011????0??????01: c_nzimm18hi = '1;
32'b????????????????011???1???????01: c_nzimm18hi = '1;
32'b????????????????011?1?????????01: c_nzimm18hi = '1;
32'b????????????????011?????1?????01: c_nzimm18hi = '1;
32'b????????????????011??1????????01: c_nzimm18hi = '1;
32'b????????????????011????0??????01: c_nzimm18hi = '1;
32'b????????????????011???1???????01: c_nzimm18hi = '1;
32'b????????????????011?1?????????01: c_nzimm18hi = '1;
32'b????????????????011?????1?????01: c_nzimm18hi = '1;
32'b????????????????011??1????????01: c_nzimm18hi = '1;
32'b????????????????011????0??????01: c_nzimm18hi = '1;
32'b????????????????011???1???????01: c_nzimm18hi = '1;
32'b????????????????011?1?????????01: c_nzimm18hi = '1;
32'b????????????????011?????1?????01: c_nzimm18hi = '1;
32'b????????????????011??1????????01: c_nzimm18hi = '1;
32'b????????????????011????0??????01: c_nzimm18hi = '1;
32'b????????????????011???1???????01: c_nzimm18hi = '1;
32'b????????????????011?1?????????01: c_nzimm18hi = '1;
32'b????????????????011?????1?????01: c_nzimm18hi = '1;
32'b????????????????011??1????????01: c_nzimm18hi = '1;
32'b????????????????011????0??????01: c_nzimm18hi = '1;
32'b????????????????011???1???????01: c_nzimm18hi = '1;
default: c_nzimm18hi = '0;
endcase
return c_nzimm18hi;
endfunction
function automatic logic riscv_decode_c_nzimm18lo(
input logic [31:0] data
);
logic c_nzimm18lo;
casez (data[31:0])
32'b????????????????011?1?????????01: c_nzimm18lo = '1;
32'b????????????????011?????1?????01: c_nzimm18lo = '1;
32'b????????????????011??1????????01: c_nzimm18lo = '1;
32'b????????????????011????0??????01: c_nzimm18lo = '1;
32'b????????????????011???1???????01: c_nzimm18lo = '1;
32'b????????????????011?1?????????01: c_nzimm18lo = '1;
32'b????????????????011?????1?????01: c_nzimm18lo = '1;
32'b????????????????011??1????????01: c_nzimm18lo = '1;
32'b????????????????011????0??????01: c_nzimm18lo = '1;
32'b????????????????011???1???????01: c_nzimm18lo = '1;
32'b????????????????011?1?????????01: c_nzimm18lo = '1;
32'b????????????????011?????1?????01: c_nzimm18lo = '1;
32'b????????????????011??1????????01: c_nzimm18lo = '1;
32'b????????????????011????0??????01: c_nzimm18lo = '1;
32'b????????????????011???1???????01: c_nzimm18lo = '1;
32'b????????????????011?1?????????01: c_nzimm18lo = '1;
32'b????????????????011?????1?????01: c_nzimm18lo = '1;
32'b????????????????011??1????????01: c_nzimm18lo = '1;
32'b????????????????011????0??????01: c_nzimm18lo = '1;
32'b????????????????011???1???????01: c_nzimm18lo = '1;
32'b????????????????011?1?????????01: c_nzimm18lo = '1;
32'b????????????????011?????1?????01: c_nzimm18lo = '1;
32'b????????????????011??1????????01: c_nzimm18lo = '1;
32'b????????????????011????0??????01: c_nzimm18lo = '1;
32'b????????????????011???1???????01: c_nzimm18lo = '1;
default: c_nzimm18lo = '0;
endcase
return c_nzimm18lo;
endfunction
function automatic logic riscv_decode_c_nzimm6hi(
input logic [31:0] data
);
logic c_nzimm6hi;
casez (data[31:0])
32'b????????????????000?1?????????01: c_nzimm6hi = '1;
32'b????????????????000??1????????01: c_nzimm6hi = '1;
32'b????????????????000?????1?????01: c_nzimm6hi = '1;
32'b????????????????000???1???????01: c_nzimm6hi = '1;
32'b????????????????000????1??????01: c_nzimm6hi = '1;
32'b????????????????000?1?????????01: c_nzimm6hi = '1;
32'b????????????????000??1????????01: c_nzimm6hi = '1;
32'b????????????????000?????1?????01: c_nzimm6hi = '1;
32'b????????????????000???1???????01: c_nzimm6hi = '1;
32'b????????????????000????1??????01: c_nzimm6hi = '1;
32'b????????????????000?1?????????01: c_nzimm6hi = '1;
32'b????????????????000??1????????01: c_nzimm6hi = '1;
32'b????????????????000?????1?????01: c_nzimm6hi = '1;
32'b????????????????000???1???????01: c_nzimm6hi = '1;
32'b????????????????000????1??????01: c_nzimm6hi = '1;
32'b????????????????000?1?????????01: c_nzimm6hi = '1;
32'b????????????????000??1????????01: c_nzimm6hi = '1;
32'b????????????????000?????1?????01: c_nzimm6hi = '1;
32'b????????????????000???1???????01: c_nzimm6hi = '1;
32'b????????????????000????1??????01: c_nzimm6hi = '1;
32'b????????????????000?1?????????01: c_nzimm6hi = '1;
32'b????????????????000??1????????01: c_nzimm6hi = '1;
32'b????????????????000?????1?????01: c_nzimm6hi = '1;
32'b????????????????000???1???????01: c_nzimm6hi = '1;
32'b????????????????000????1??????01: c_nzimm6hi = '1;
32'b????????????????000?00000?????01: c_nzimm6hi = '1;
default: c_nzimm6hi = '0;
endcase
return c_nzimm6hi;
endfunction
function automatic logic riscv_decode_c_nzimm6lo(
input logic [31:0] data
);
logic c_nzimm6lo;
casez (data[31:0])
32'b????????????????000?1?????????01: c_nzimm6lo = '1;
32'b????????????????000??1????????01: c_nzimm6lo = '1;
32'b????????????????000?????1?????01: c_nzimm6lo = '1;
32'b????????????????000???1???????01: c_nzimm6lo = '1;
32'b????????????????000????1??????01: c_nzimm6lo = '1;
32'b????????????????000?1?????????01: c_nzimm6lo = '1;
32'b????????????????000??1????????01: c_nzimm6lo = '1;
32'b????????????????000?????1?????01: c_nzimm6lo = '1;
32'b????????????????000???1???????01: c_nzimm6lo = '1;
32'b????????????????000????1??????01: c_nzimm6lo = '1;
32'b????????????????000?1?????????01: c_nzimm6lo = '1;
32'b????????????????000??1????????01: c_nzimm6lo = '1;
32'b????????????????000?????1?????01: c_nzimm6lo = '1;
32'b????????????????000???1???????01: c_nzimm6lo = '1;
32'b????????????????000????1??????01: c_nzimm6lo = '1;
32'b????????????????000?1?????????01: c_nzimm6lo = '1;
32'b????????????????000??1????????01: c_nzimm6lo = '1;
32'b????????????????000?????1?????01: c_nzimm6lo = '1;
32'b????????????????000???1???????01: c_nzimm6lo = '1;
32'b????????????????000????1??????01: c_nzimm6lo = '1;
32'b????????????????000?1?????????01: c_nzimm6lo = '1;
32'b????????????????000??1????????01: c_nzimm6lo = '1;
32'b????????????????000?????1?????01: c_nzimm6lo = '1;
32'b????????????????000???1???????01: c_nzimm6lo = '1;
32'b????????????????000????1??????01: c_nzimm6lo = '1;
32'b????????????????000?00000?????01: c_nzimm6lo = '1;
default: c_nzimm6lo = '0;
endcase
return c_nzimm6lo;
endfunction
function automatic logic riscv_decode_c_nzuimm10(
input logic [31:0] data
);
logic c_nzuimm10;
casez (data[31:0])
32'b????????????????000???????????00: c_nzuimm10 = '1;
default: c_nzuimm10 = '0;
endcase
return c_nzuimm10;
endfunction
function automatic logic riscv_decode_c_nzuimm6hi(
input logic [31:0] data
);
logic c_nzuimm6hi;
casez (data[31:0])
32'b????????????????000???1???????10: c_nzuimm6hi = '1;
32'b????????????????000?????1?????10: c_nzuimm6hi = '1;
32'b????????????????000????1??????10: c_nzuimm6hi = '1;
32'b????????????????000?1?????????10: c_nzuimm6hi = '1;
32'b????????????????000??1????????10: c_nzuimm6hi = '1;
32'b????????????????000???1???????10: c_nzuimm6hi = '1;
32'b????????????????000?????1?????10: c_nzuimm6hi = '1;
32'b????????????????000????1??????10: c_nzuimm6hi = '1;
32'b????????????????000?1?????????10: c_nzuimm6hi = '1;
32'b????????????????000??1????????10: c_nzuimm6hi = '1;
32'b????????????????000???1???????10: c_nzuimm6hi = '1;
32'b????????????????000?????1?????10: c_nzuimm6hi = '1;
32'b????????????????000????1??????10: c_nzuimm6hi = '1;
32'b????????????????000?1?????????10: c_nzuimm6hi = '1;
32'b????????????????000??1????????10: c_nzuimm6hi = '1;
32'b????????????????000???1???????10: c_nzuimm6hi = '1;
32'b????????????????000?????1?????10: c_nzuimm6hi = '1;
32'b????????????????000????1??????10: c_nzuimm6hi = '1;
32'b????????????????000?1?????????10: c_nzuimm6hi = '1;
32'b????????????????000??1????????10: c_nzuimm6hi = '1;
32'b????????????????000???1???????10: c_nzuimm6hi = '1;
32'b????????????????000?????1?????10: c_nzuimm6hi = '1;
32'b????????????????000????1??????10: c_nzuimm6hi = '1;
32'b????????????????000?1?????????10: c_nzuimm6hi = '1;
32'b????????????????000??1????????10: c_nzuimm6hi = '1;
32'b????????????????100?01????????01: c_nzuimm6hi = '1;
32'b????????????????100?00????????01: c_nzuimm6hi = '1;
default: c_nzuimm6hi = '0;
endcase
return c_nzuimm6hi;
endfunction
function automatic logic riscv_decode_c_nzuimm6lo(
input logic [31:0] data
);
logic c_nzuimm6lo;
casez (data[31:0])
32'b????????????????000???1???????10: c_nzuimm6lo = '1;
32'b????????????????000?????1?????10: c_nzuimm6lo = '1;
32'b????????????????000????1??????10: c_nzuimm6lo = '1;
32'b????????????????000?1?????????10: c_nzuimm6lo = '1;
32'b????????????????000??1????????10: c_nzuimm6lo = '1;
32'b????????????????000???1???????10: c_nzuimm6lo = '1;
32'b????????????????000?????1?????10: c_nzuimm6lo = '1;
32'b????????????????000????1??????10: c_nzuimm6lo = '1;
32'b????????????????000?1?????????10: c_nzuimm6lo = '1;
32'b????????????????000??1????????10: c_nzuimm6lo = '1;
32'b????????????????000???1???????10: c_nzuimm6lo = '1;
32'b????????????????000?????1?????10: c_nzuimm6lo = '1;
32'b????????????????000????1??????10: c_nzuimm6lo = '1;
32'b????????????????000?1?????????10: c_nzuimm6lo = '1;
32'b????????????????000??1????????10: c_nzuimm6lo = '1;
32'b????????????????000???1???????10: c_nzuimm6lo = '1;
32'b????????????????000?????1?????10: c_nzuimm6lo = '1;
32'b????????????????000????1??????10: c_nzuimm6lo = '1;
32'b????????????????000?1?????????10: c_nzuimm6lo = '1;
32'b????????????????000??1????????10: c_nzuimm6lo = '1;
32'b????????????????000???1???????10: c_nzuimm6lo = '1;
32'b????????????????000?????1?????10: c_nzuimm6lo = '1;
32'b????????????????000????1??????10: c_nzuimm6lo = '1;
32'b????????????????000?1?????????10: c_nzuimm6lo = '1;
32'b????????????????000??1????????10: c_nzuimm6lo = '1;
32'b????????????????100?01????????01: c_nzuimm6lo = '1;
32'b????????????????100?00????????01: c_nzuimm6lo = '1;
default: c_nzuimm6lo = '0;
endcase
return c_nzuimm6lo;
endfunction
function automatic logic riscv_decode_c_rs2(
input logic [31:0] data
);
logic c_rs2;
casez (data[31:0])
32'b????????????????1001????????1?10: c_rs2 = '1;
32'b????????????????1001??????1???10: c_rs2 = '1;
32'b????????????????1001???????1??10: c_rs2 = '1;
32'b????????????????1001?????1????10: c_rs2 = '1;
32'b????????????????1001?????????110: c_rs2 = '1;
32'b????????????????1001????????1?10: c_rs2 = '1;
32'b????????????????1001??????1???10: c_rs2 = '1;
32'b????????????????1001???????1??10: c_rs2 = '1;
32'b????????????????1001?????1????10: c_rs2 = '1;
32'b????????????????1001?????????110: c_rs2 = '1;
32'b????????????????1001????????1?10: c_rs2 = '1;
32'b????????????????1001??????1???10: c_rs2 = '1;
32'b????????????????1001???????1??10: c_rs2 = '1;
32'b????????????????1001?????1????10: c_rs2 = '1;
32'b????????????????1001?????????110: c_rs2 = '1;
32'b????????????????1001????????1?10: c_rs2 = '1;
32'b????????????????1001??????1???10: c_rs2 = '1;
32'b????????????????1001???????1??10: c_rs2 = '1;
32'b????????????????1001?????1????10: c_rs2 = '1;
32'b????????????????1001?????????110: c_rs2 = '1;
32'b????????????????1001????????1?10: c_rs2 = '1;
32'b????????????????1001??????1???10: c_rs2 = '1;
32'b????????????????1001???????1??10: c_rs2 = '1;
32'b????????????????1001?????1????10: c_rs2 = '1;
32'b????????????????1001?????????110: c_rs2 = '1;
32'b????????????????1000?????1????10: c_rs2 = '1;
32'b????????????????1000???????1??10: c_rs2 = '1;
32'b????????????????1000?????????110: c_rs2 = '1;
32'b????????????????1000????????1?10: c_rs2 = '1;
32'b????????????????1000??????1???10: c_rs2 = '1;
32'b????????????????1000?????1????10: c_rs2 = '1;
32'b????????????????1000???????1??10: c_rs2 = '1;
32'b????????????????1000?????????110: c_rs2 = '1;
32'b????????????????1000????????1?10: c_rs2 = '1;
32'b????????????????1000??????1???10: c_rs2 = '1;
32'b????????????????1000?????1????10: c_rs2 = '1;
32'b????????????????1000???????1??10: c_rs2 = '1;
32'b????????????????1000?????????110: c_rs2 = '1;
32'b????????????????1000????????1?10: c_rs2 = '1;
32'b????????????????1000??????1???10: c_rs2 = '1;
32'b????????????????1000?????1????10: c_rs2 = '1;
32'b????????????????1000???????1??10: c_rs2 = '1;
32'b????????????????1000?????????110: c_rs2 = '1;
32'b????????????????1000????????1?10: c_rs2 = '1;
32'b????????????????1000??????1???10: c_rs2 = '1;
32'b????????????????1000?????1????10: c_rs2 = '1;
32'b????????????????1000???????1??10: c_rs2 = '1;
32'b????????????????1000?????????110: c_rs2 = '1;
32'b????????????????1000????????1?10: c_rs2 = '1;
32'b????????????????1000??????1???10: c_rs2 = '1;
32'b????????????????110???????????10: c_rs2 = '1;
default: c_rs2 = '0;
endcase
return c_rs2;
endfunction
function automatic logic riscv_decode_c_uimm7hi(
input logic [31:0] data
);
logic c_uimm7hi;
casez (data[31:0])
32'b????????????????010???????????00: c_uimm7hi = '1;
32'b????????????????110???????????00: c_uimm7hi = '1;
default: c_uimm7hi = '0;
endcase
return c_uimm7hi;
endfunction
function automatic logic riscv_decode_c_uimm7lo(
input logic [31:0] data
);
logic c_uimm7lo;
casez (data[31:0])
32'b????????????????010???????????00: c_uimm7lo = '1;
32'b????????????????110???????????00: c_uimm7lo = '1;
default: c_uimm7lo = '0;
endcase
return c_uimm7lo;
endfunction
function automatic logic riscv_decode_c_uimm8sp_s(
input logic [31:0] data
);
logic c_uimm8sp_s;
casez (data[31:0])
32'b????????????????110???????????10: c_uimm8sp_s = '1;
default: c_uimm8sp_s = '0;
endcase
return c_uimm8sp_s;
endfunction
function automatic logic riscv_decode_c_uimm8sphi(
input logic [31:0] data
);
logic c_uimm8sphi;
casez (data[31:0])
32'b????????????????010????1??????10: c_uimm8sphi = '1;
32'b????????????????010???1???????10: c_uimm8sphi = '1;
32'b????????????????010??1????????10: c_uimm8sphi = '1;
32'b????????????????010?1?????????10: c_uimm8sphi = '1;
32'b????????????????010?????1?????10: c_uimm8sphi = '1;
32'b????????????????010????1??????10: c_uimm8sphi = '1;
32'b????????????????010???1???????10: c_uimm8sphi = '1;
32'b????????????????010??1????????10: c_uimm8sphi = '1;
32'b????????????????010?1?????????10: c_uimm8sphi = '1;
32'b????????????????010?????1?????10: c_uimm8sphi = '1;
32'b????????????????010????1??????10: c_uimm8sphi = '1;
32'b????????????????010???1???????10: c_uimm8sphi = '1;
32'b????????????????010??1????????10: c_uimm8sphi = '1;
32'b????????????????010?1?????????10: c_uimm8sphi = '1;
32'b????????????????010?????1?????10: c_uimm8sphi = '1;
32'b????????????????010????1??????10: c_uimm8sphi = '1;
32'b????????????????010???1???????10: c_uimm8sphi = '1;
32'b????????????????010??1????????10: c_uimm8sphi = '1;
32'b????????????????010?1?????????10: c_uimm8sphi = '1;
32'b????????????????010?????1?????10: c_uimm8sphi = '1;
32'b????????????????010????1??????10: c_uimm8sphi = '1;
32'b????????????????010???1???????10: c_uimm8sphi = '1;
32'b????????????????010??1????????10: c_uimm8sphi = '1;
32'b????????????????010?1?????????10: c_uimm8sphi = '1;
32'b????????????????010?????1?????10: c_uimm8sphi = '1;
default: c_uimm8sphi = '0;
endcase
return c_uimm8sphi;
endfunction
function automatic logic riscv_decode_c_uimm8splo(
input logic [31:0] data
);
logic c_uimm8splo;
casez (data[31:0])
32'b????????????????010????1??????10: c_uimm8splo = '1;
32'b????????????????010???1???????10: c_uimm8splo = '1;
32'b????????????????010??1????????10: c_uimm8splo = '1;
32'b????????????????010?1?????????10: c_uimm8splo = '1;
32'b????????????????010?????1?????10: c_uimm8splo = '1;
32'b????????????????010????1??????10: c_uimm8splo = '1;
32'b????????????????010???1???????10: c_uimm8splo = '1;
32'b????????????????010??1????????10: c_uimm8splo = '1;
32'b????????????????010?1?????????10: c_uimm8splo = '1;
32'b????????????????010?????1?????10: c_uimm8splo = '1;
32'b????????????????010????1??????10: c_uimm8splo = '1;
32'b????????????????010???1???????10: c_uimm8splo = '1;
32'b????????????????010??1????????10: c_uimm8splo = '1;
32'b????????????????010?1?????????10: c_uimm8splo = '1;
32'b????????????????010?????1?????10: c_uimm8splo = '1;
32'b????????????????010????1??????10: c_uimm8splo = '1;
32'b????????????????010???1???????10: c_uimm8splo = '1;
32'b????????????????010??1????????10: c_uimm8splo = '1;
32'b????????????????010?1?????????10: c_uimm8splo = '1;
32'b????????????????010?????1?????10: c_uimm8splo = '1;
32'b????????????????010????1??????10: c_uimm8splo = '1;
32'b????????????????010???1???????10: c_uimm8splo = '1;
32'b????????????????010??1????????10: c_uimm8splo = '1;
32'b????????????????010?1?????????10: c_uimm8splo = '1;
32'b????????????????010?????1?????10: c_uimm8splo = '1;
default: c_uimm8splo = '0;
endcase
return c_uimm8splo;
endfunction
function automatic logic riscv_decode_fm(
input logic [31:0] data
);
logic fm;
casez (data[31:0])
32'b?????????????????000?????0001111: fm = '1;
default: fm = '0;
endcase
return fm;
endfunction
function automatic logic riscv_decode_imm12(
input logic [31:0] data
);
logic imm12;
casez (data[31:0])
32'b?????????????????000?????0010011: imm12 = '1;
32'b?????????????????111?????0010011: imm12 = '1;
32'b?????????????????000?????1100111: imm12 = '1;
32'b?????????????????000?????0000011: imm12 = '1;
32'b?????????????????100?????0000011: imm12 = '1;
32'b?????????????????001?????0000011: imm12 = '1;
32'b?????????????????101?????0000011: imm12 = '1;
32'b?????????????????010?????0000011: imm12 = '1;
32'b?????????????????110?????0010011: imm12 = '1;
32'b?????????????????010?????0010011: imm12 = '1;
32'b?????????????????011?????0010011: imm12 = '1;
32'b?????????????????100?????0010011: imm12 = '1;
default: imm12 = '0;
endcase
return imm12;
endfunction
function automatic logic riscv_decode_imm12hi(
input logic [31:0] data
);
logic imm12hi;
casez (data[31:0])
32'b?????????????????000?????0100011: imm12hi = '1;
32'b?????????????????001?????0100011: imm12hi = '1;
32'b?????????????????010?????0100011: imm12hi = '1;
default: imm12hi = '0;
endcase
return imm12hi;
endfunction
function automatic logic riscv_decode_imm12lo(
input logic [31:0] data
);
logic imm12lo;
casez (data[31:0])
32'b?????????????????000?????0100011: imm12lo = '1;
32'b?????????????????001?????0100011: imm12lo = '1;
32'b?????????????????010?????0100011: imm12lo = '1;
default: imm12lo = '0;
endcase
return imm12lo;
endfunction
function automatic logic riscv_decode_imm20(
input logic [31:0] data
);
logic imm20;
casez (data[31:0])
32'b?????????????????????????0010111: imm20 = '1;
32'b?????????????????????????0110111: imm20 = '1;
default: imm20 = '0;
endcase
return imm20;
endfunction
function automatic logic riscv_decode_jimm20(
input logic [31:0] data
);
logic jimm20;
casez (data[31:0])
32'b?????????????????????????1101111: jimm20 = '1;
default: jimm20 = '0;
endcase
return jimm20;
endfunction
function automatic logic riscv_decode_pred(
input logic [31:0] data
);
logic pred;
casez (data[31:0])
32'b?????????????????000?????0001111: pred = '1;
default: pred = '0;
endcase
return pred;
endfunction
function automatic logic riscv_decode_rd(
input logic [31:0] data
);
logic rd;
casez (data[31:0])
32'b0000000??????????000?????0110011: rd = '1;
32'b?????????????????000?????0010011: rd = '1;
32'b0000000??????????111?????0110011: rd = '1;
32'b?????????????????111?????0010011: rd = '1;
32'b?????????????????????????0010111: rd = '1;
32'b????????????????010???????????01: rd = '1;
32'b????????????????011?1?????????01: rd = '1;
32'b????????????????011?????1?????01: rd = '1;
32'b????????????????011??1????????01: rd = '1;
32'b????????????????011????0??????01: rd = '1;
32'b????????????????011???1???????01: rd = '1;
32'b????????????????011?1?????????01: rd = '1;
32'b????????????????011?????1?????01: rd = '1;
32'b????????????????011??1????????01: rd = '1;
32'b????????????????011????0??????01: rd = '1;
32'b????????????????011???1???????01: rd = '1;
32'b????????????????011?1?????????01: rd = '1;
32'b????????????????011?????1?????01: rd = '1;
32'b????????????????011??1????????01: rd = '1;
32'b????????????????011????0??????01: rd = '1;
32'b????????????????011???1???????01: rd = '1;
32'b????????????????011?1?????????01: rd = '1;
32'b????????????????011?????1?????01: rd = '1;
32'b????????????????011??1????????01: rd = '1;
32'b????????????????011????0??????01: rd = '1;
32'b????????????????011???1???????01: rd = '1;
32'b????????????????011?1?????????01: rd = '1;
32'b????????????????011?????1?????01: rd = '1;
32'b????????????????011??1????????01: rd = '1;
32'b????????????????011????0??????01: rd = '1;
32'b????????????????011???1???????01: rd = '1;
32'b????????????????010????1??????10: rd = '1;
32'b????????????????010???1???????10: rd = '1;
32'b????????????????010??1????????10: rd = '1;
32'b????????????????010?1?????????10: rd = '1;
32'b????????????????010?????1?????10: rd = '1;
32'b????????????????010????1??????10: rd = '1;
32'b????????????????010???1???????10: rd = '1;
32'b????????????????010??1????????10: rd = '1;
32'b????????????????010?1?????????10: rd = '1;
32'b????????????????010?????1?????10: rd = '1;
32'b????????????????010????1??????10: rd = '1;
32'b????????????????010???1???????10: rd = '1;
32'b????????????????010??1????????10: rd = '1;
32'b????????????????010?1?????????10: rd = '1;
32'b????????????????010?????1?????10: rd = '1;
32'b????????????????010????1??????10: rd = '1;
32'b????????????????010???1???????10: rd = '1;
32'b????????????????010??1????????10: rd = '1;
32'b????????????????010?1?????????10: rd = '1;
32'b????????????????010?????1?????10: rd = '1;
32'b????????????????010????1??????10: rd = '1;
32'b????????????????010???1???????10: rd = '1;
32'b????????????????010??1????????10: rd = '1;
32'b????????????????010?1?????????10: rd = '1;
32'b????????????????010?????1?????10: rd = '1;
32'b????????????????1000?????1????10: rd = '1;
32'b????????????????1000???????1??10: rd = '1;
32'b????????????????1000?????????110: rd = '1;
32'b????????????????1000????????1?10: rd = '1;
32'b????????????????1000??????1???10: rd = '1;
32'b????????????????1000?????1????10: rd = '1;
32'b????????????????1000???????1??10: rd = '1;
32'b????????????????1000?????????110: rd = '1;
32'b????????????????1000????????1?10: rd = '1;
32'b????????????????1000??????1???10: rd = '1;
32'b????????????????1000?????1????10: rd = '1;
32'b????????????????1000???????1??10: rd = '1;
32'b????????????????1000?????????110: rd = '1;
32'b????????????????1000????????1?10: rd = '1;
32'b????????????????1000??????1???10: rd = '1;
32'b????????????????1000?????1????10: rd = '1;
32'b????????????????1000???????1??10: rd = '1;
32'b????????????????1000?????????110: rd = '1;
32'b????????????????1000????????1?10: rd = '1;
32'b????????????????1000??????1???10: rd = '1;
32'b????????????????1000?????1????10: rd = '1;
32'b????????????????1000???????1??10: rd = '1;
32'b????????????????1000?????????110: rd = '1;
32'b????????????????1000????????1?10: rd = '1;
32'b????????????????1000??????1???10: rd = '1;
32'b0000001??????????100?????0110011: rd = '1;
32'b0000001??????????101?????0110011: rd = '1;
32'b?????????????????000?????0001111: rd = '1;
32'b?????????????????????????1101111: rd = '1;
32'b?????????????????000?????1100111: rd = '1;
32'b?????????????????000?????0000011: rd = '1;
32'b?????????????????100?????0000011: rd = '1;
32'b?????????????????001?????0000011: rd = '1;
32'b?????????????????101?????0000011: rd = '1;
32'b?????????????????????????0110111: rd = '1;
32'b?????????????????010?????0000011: rd = '1;
32'b0000001??????????000?????0110011: rd = '1;
32'b0000001??????????001?????0110011: rd = '1;
32'b0000001??????????010?????0110011: rd = '1;
32'b0000001??????????011?????0110011: rd = '1;
32'b0000000??????????110?????0110011: rd = '1;
32'b?????????????????110?????0010011: rd = '1;
32'b0000001??????????110?????0110011: rd = '1;
32'b0000001??????????111?????0110011: rd = '1;
32'b0000000??????????001?????0110011: rd = '1;
32'b000000???????????001?????0010011: rd = '1;
32'b0000000??????????010?????0110011: rd = '1;
32'b?????????????????010?????0010011: rd = '1;
32'b?????????????????011?????0010011: rd = '1;
32'b0000000??????????011?????0110011: rd = '1;
32'b0100000??????????101?????0110011: rd = '1;
32'b010000???????????101?????0010011: rd = '1;
32'b0000000??????????101?????0110011: rd = '1;
32'b000000???????????101?????0010011: rd = '1;
32'b0100000??????????000?????0110011: rd = '1;
32'b0000000??????????100?????0110011: rd = '1;
32'b?????????????????100?????0010011: rd = '1;
default: rd = '0;
endcase
return rd;
endfunction
function automatic logic riscv_decode_rd_p(
input logic [31:0] data
);
logic rd_p;
casez (data[31:0])
32'b????????????????000???????????00: rd_p = '1;
32'b????????????????010???????????00: rd_p = '1;
default: rd_p = '0;
endcase
return rd_p;
endfunction
function automatic logic riscv_decode_rd_rs1(
input logic [31:0] data
);
logic rd_rs1;
casez (data[31:0])
32'b????????????????1001????????1?10: rd_rs1 = '1;
32'b????????????????1001??????1???10: rd_rs1 = '1;
32'b????????????????1001???????1??10: rd_rs1 = '1;
32'b????????????????1001?????1????10: rd_rs1 = '1;
32'b????????????????1001?????????110: rd_rs1 = '1;
32'b????????????????1001????????1?10: rd_rs1 = '1;
32'b????????????????1001??????1???10: rd_rs1 = '1;
32'b????????????????1001???????1??10: rd_rs1 = '1;
32'b????????????????1001?????1????10: rd_rs1 = '1;
32'b????????????????1001?????????110: rd_rs1 = '1;
32'b????????????????1001????????1?10: rd_rs1 = '1;
32'b????????????????1001??????1???10: rd_rs1 = '1;
32'b????????????????1001???????1??10: rd_rs1 = '1;
32'b????????????????1001?????1????10: rd_rs1 = '1;
32'b????????????????1001?????????110: rd_rs1 = '1;
32'b????????????????1001????????1?10: rd_rs1 = '1;
32'b????????????????1001??????1???10: rd_rs1 = '1;
32'b????????????????1001???????1??10: rd_rs1 = '1;
32'b????????????????1001?????1????10: rd_rs1 = '1;
32'b????????????????1001?????????110: rd_rs1 = '1;
32'b????????????????1001????????1?10: rd_rs1 = '1;
32'b????????????????1001??????1???10: rd_rs1 = '1;
32'b????????????????1001???????1??10: rd_rs1 = '1;
32'b????????????????1001?????1????10: rd_rs1 = '1;
32'b????????????????1001?????????110: rd_rs1 = '1;
32'b????????????????000?1?????????01: rd_rs1 = '1;
32'b????????????????000??1????????01: rd_rs1 = '1;
32'b????????????????000?????1?????01: rd_rs1 = '1;
32'b????????????????000???1???????01: rd_rs1 = '1;
32'b????????????????000????1??????01: rd_rs1 = '1;
32'b????????????????000?1?????????01: rd_rs1 = '1;
32'b????????????????000??1????????01: rd_rs1 = '1;
32'b????????????????000?????1?????01: rd_rs1 = '1;
32'b????????????????000???1???????01: rd_rs1 = '1;
32'b????????????????000????1??????01: rd_rs1 = '1;
32'b????????????????000?1?????????01: rd_rs1 = '1;
32'b????????????????000??1????????01: rd_rs1 = '1;
32'b????????????????000?????1?????01: rd_rs1 = '1;
32'b????????????????000???1???????01: rd_rs1 = '1;
32'b????????????????000????1??????01: rd_rs1 = '1;
32'b????????????????000?1?????????01: rd_rs1 = '1;
32'b????????????????000??1????????01: rd_rs1 = '1;
32'b????????????????000?????1?????01: rd_rs1 = '1;
32'b????????????????000???1???????01: rd_rs1 = '1;
32'b????????????????000????1??????01: rd_rs1 = '1;
32'b????????????????000?1?????????01: rd_rs1 = '1;
32'b????????????????000??1????????01: rd_rs1 = '1;
32'b????????????????000?????1?????01: rd_rs1 = '1;
32'b????????????????000???1???????01: rd_rs1 = '1;
32'b????????????????000????1??????01: rd_rs1 = '1;
32'b????????????????000???1???????10: rd_rs1 = '1;
32'b????????????????000?????1?????10: rd_rs1 = '1;
32'b????????????????000????1??????10: rd_rs1 = '1;
32'b????????????????000?1?????????10: rd_rs1 = '1;
32'b????????????????000??1????????10: rd_rs1 = '1;
32'b????????????????000???1???????10: rd_rs1 = '1;
32'b????????????????000?????1?????10: rd_rs1 = '1;
32'b????????????????000????1??????10: rd_rs1 = '1;
32'b????????????????000?1?????????10: rd_rs1 = '1;
32'b????????????????000??1????????10: rd_rs1 = '1;
32'b????????????????000???1???????10: rd_rs1 = '1;
32'b????????????????000?????1?????10: rd_rs1 = '1;
32'b????????????????000????1??????10: rd_rs1 = '1;
32'b????????????????000?1?????????10: rd_rs1 = '1;
32'b????????????????000??1????????10: rd_rs1 = '1;
32'b????????????????000???1???????10: rd_rs1 = '1;
32'b????????????????000?????1?????10: rd_rs1 = '1;
32'b????????????????000????1??????10: rd_rs1 = '1;
32'b????????????????000?1?????????10: rd_rs1 = '1;
32'b????????????????000??1????????10: rd_rs1 = '1;
32'b????????????????000???1???????10: rd_rs1 = '1;
32'b????????????????000?????1?????10: rd_rs1 = '1;
32'b????????????????000????1??????10: rd_rs1 = '1;
32'b????????????????000?1?????????10: rd_rs1 = '1;
32'b????????????????000??1????????10: rd_rs1 = '1;
default: rd_rs1 = '0;
endcase
return rd_rs1;
endfunction
function automatic logic riscv_decode_rd_rs1_p(
input logic [31:0] data
);
logic rd_rs1_p;
casez (data[31:0])
32'b????????????????100011???11???01: rd_rs1_p = '1;
32'b????????????????100?10????????01: rd_rs1_p = '1;
32'b????????????????100011???10???01: rd_rs1_p = '1;
32'b????????????????100?01????????01: rd_rs1_p = '1;
32'b????????????????100?00????????01: rd_rs1_p = '1;
32'b????????????????100011???00???01: rd_rs1_p = '1;
32'b????????????????100011???01???01: rd_rs1_p = '1;
default: rd_rs1_p = '0;
endcase
return rd_rs1_p;
endfunction
function automatic logic riscv_decode_rs1(
input logic [31:0] data
);
logic rs1;
casez (data[31:0])
32'b0000000??????????000?????0110011: rs1 = '1;
32'b?????????????????000?????0010011: rs1 = '1;
32'b0000000??????????111?????0110011: rs1 = '1;
32'b?????????????????111?????0010011: rs1 = '1;
32'b?????????????????000?????1100011: rs1 = '1;
32'b?????????????????101?????1100011: rs1 = '1;
32'b?????????????????111?????1100011: rs1 = '1;
32'b?????????????????100?????1100011: rs1 = '1;
32'b?????????????????110?????1100011: rs1 = '1;
32'b?????????????????001?????1100011: rs1 = '1;
32'b????????????????1000?????0000010: rs1 = '1;
32'b0000001??????????100?????0110011: rs1 = '1;
32'b0000001??????????101?????0110011: rs1 = '1;
32'b?????????????????000?????0001111: rs1 = '1;
32'b?????????????????000?????1100111: rs1 = '1;
32'b?????????????????000?????0000011: rs1 = '1;
32'b?????????????????100?????0000011: rs1 = '1;
32'b?????????????????001?????0000011: rs1 = '1;
32'b?????????????????101?????0000011: rs1 = '1;
32'b?????????????????010?????0000011: rs1 = '1;
32'b0000001??????????000?????0110011: rs1 = '1;
32'b0000001??????????001?????0110011: rs1 = '1;
32'b0000001??????????010?????0110011: rs1 = '1;
32'b0000001??????????011?????0110011: rs1 = '1;
32'b0000000??????????110?????0110011: rs1 = '1;
32'b?????????????????110?????0010011: rs1 = '1;
32'b0000001??????????110?????0110011: rs1 = '1;
32'b0000001??????????111?????0110011: rs1 = '1;
32'b?????????????????000?????0100011: rs1 = '1;
32'b?????????????????001?????0100011: rs1 = '1;
32'b0000000??????????001?????0110011: rs1 = '1;
32'b000000???????????001?????0010011: rs1 = '1;
32'b0000000??????????010?????0110011: rs1 = '1;
32'b?????????????????010?????0010011: rs1 = '1;
32'b?????????????????011?????0010011: rs1 = '1;
32'b0000000??????????011?????0110011: rs1 = '1;
32'b0100000??????????101?????0110011: rs1 = '1;
32'b010000???????????101?????0010011: rs1 = '1;
32'b0000000??????????101?????0110011: rs1 = '1;
32'b000000???????????101?????0010011: rs1 = '1;
32'b0100000??????????000?????0110011: rs1 = '1;
32'b?????????????????010?????0100011: rs1 = '1;
32'b0000000??????????100?????0110011: rs1 = '1;
32'b?????????????????100?????0010011: rs1 = '1;
default: rs1 = '0;
endcase
return rs1;
endfunction
function automatic logic riscv_decode_rs1_p(
input logic [31:0] data
);
logic rs1_p;
casez (data[31:0])
32'b????????????????110???????????01: rs1_p = '1;
32'b????????????????111???????????01: rs1_p = '1;
32'b????????????????010???????????00: rs1_p = '1;
32'b????????????????110???????????00: rs1_p = '1;
default: rs1_p = '0;
endcase
return rs1_p;
endfunction
function automatic logic riscv_decode_rs2(
input logic [31:0] data
);
logic rs2;
casez (data[31:0])
32'b0000000??????????000?????0110011: rs2 = '1;
32'b0000000??????????111?????0110011: rs2 = '1;
32'b?????????????????000?????1100011: rs2 = '1;
32'b?????????????????101?????1100011: rs2 = '1;
32'b?????????????????111?????1100011: rs2 = '1;
32'b?????????????????100?????1100011: rs2 = '1;
32'b?????????????????110?????1100011: rs2 = '1;
32'b?????????????????001?????1100011: rs2 = '1;
32'b0000001??????????100?????0110011: rs2 = '1;
32'b0000001??????????101?????0110011: rs2 = '1;
32'b0000001??????????000?????0110011: rs2 = '1;
32'b0000001??????????001?????0110011: rs2 = '1;
32'b0000001??????????010?????0110011: rs2 = '1;
32'b0000001??????????011?????0110011: rs2 = '1;
32'b0000000??????????110?????0110011: rs2 = '1;
32'b0000001??????????110?????0110011: rs2 = '1;
32'b0000001??????????111?????0110011: rs2 = '1;
32'b?????????????????000?????0100011: rs2 = '1;
32'b?????????????????001?????0100011: rs2 = '1;
32'b0000000??????????001?????0110011: rs2 = '1;
32'b0000000??????????010?????0110011: rs2 = '1;
32'b0000000??????????011?????0110011: rs2 = '1;
32'b0100000??????????101?????0110011: rs2 = '1;
32'b0000000??????????101?????0110011: rs2 = '1;
32'b0100000??????????000?????0110011: rs2 = '1;
32'b?????????????????010?????0100011: rs2 = '1;
32'b0000000??????????100?????0110011: rs2 = '1;
default: rs2 = '0;
endcase
return rs2;
endfunction
function automatic logic riscv_decode_rs2_p(
input logic [31:0] data
);
logic rs2_p;
casez (data[31:0])
32'b????????????????100011???11???01: rs2_p = '1;
32'b????????????????100011???10???01: rs2_p = '1;
32'b????????????????100011???00???01: rs2_p = '1;
32'b????????????????110???????????00: rs2_p = '1;
32'b????????????????100011???01???01: rs2_p = '1;
default: rs2_p = '0;
endcase
return rs2_p;
endfunction
function automatic logic riscv_decode_shamtd(
input logic [31:0] data
);
logic shamtd;
casez (data[31:0])
32'b000000???????????001?????0010011: shamtd = '1;
32'b010000???????????101?????0010011: shamtd = '1;
32'b000000???????????101?????0010011: shamtd = '1;
default: shamtd = '0;
endcase
return shamtd;
endfunction
function automatic logic riscv_decode_succ(
input logic [31:0] data
);
logic succ;
casez (data[31:0])
32'b?????????????????000?????0001111: succ = '1;
default: succ = '0;
endcase
return succ;
endfunction
